module address_decode_6_3
(
input wire[5:0] addr_raw,
input wire selector_enabled,
output wire[63:0] addr_selector
);

wire[8:0] r_0_addr;
wire[8:0] r_1_addr;

assign r_0_addr[0] = (addr_raw[2:0]==3'b000) ?1'b1:1'b0;
assign r_0_addr[1] = (addr_raw[2:0]==3'b001) ?1'b1:1'b0;
assign r_0_addr[2] = (addr_raw[2:0]==3'b010) ?1'b1:1'b0;
assign r_0_addr[3] = (addr_raw[2:0]==3'b011) ?1'b1:1'b0;
assign r_0_addr[4] = (addr_raw[2:0]==3'b100) ?1'b1:1'b0;
assign r_0_addr[5] = (addr_raw[2:0]==3'b101) ?1'b1:1'b0;
assign r_0_addr[6] = (addr_raw[2:0]==3'b110) ?1'b1:1'b0;
assign r_0_addr[7] = (addr_raw[2:0]==3'b111) ?1'b1:1'b0;
assign r_1_addr[0] = (addr_raw[5:3]==3'b000) ?1'b1:1'b0;
assign r_1_addr[1] = (addr_raw[5:3]==3'b001) ?1'b1:1'b0;
assign r_1_addr[2] = (addr_raw[5:3]==3'b010) ?1'b1:1'b0;
assign r_1_addr[3] = (addr_raw[5:3]==3'b011) ?1'b1:1'b0;
assign r_1_addr[4] = (addr_raw[5:3]==3'b100) ?1'b1:1'b0;
assign r_1_addr[5] = (addr_raw[5:3]==3'b101) ?1'b1:1'b0;
assign r_1_addr[6] = (addr_raw[5:3]==3'b110) ?1'b1:1'b0;
assign r_1_addr[7] = (addr_raw[5:3]==3'b111) ?1'b1:1'b0;

addr_selector = {r_1_addr[7]&r_0_addr[7]&selector_enabled,
r_1_addr[7]&r_0_addr[6]&selector_enabled,
r_1_addr[7]&r_0_addr[5]&selector_enabled,
r_1_addr[7]&r_0_addr[4]&selector_enabled,
r_1_addr[7]&r_0_addr[3]&selector_enabled,
r_1_addr[7]&r_0_addr[2]&selector_enabled,
r_1_addr[7]&r_0_addr[1]&selector_enabled,
r_1_addr[7]&r_0_addr[0]&selector_enabled,
r_1_addr[6]&r_0_addr[7]&selector_enabled,
r_1_addr[6]&r_0_addr[6]&selector_enabled,
r_1_addr[6]&r_0_addr[5]&selector_enabled,
r_1_addr[6]&r_0_addr[4]&selector_enabled,
r_1_addr[6]&r_0_addr[3]&selector_enabled,
r_1_addr[6]&r_0_addr[2]&selector_enabled,
r_1_addr[6]&r_0_addr[1]&selector_enabled,
r_1_addr[6]&r_0_addr[0]&selector_enabled,
r_1_addr[5]&r_0_addr[7]&selector_enabled,
r_1_addr[5]&r_0_addr[6]&selector_enabled,
r_1_addr[5]&r_0_addr[5]&selector_enabled,
r_1_addr[5]&r_0_addr[4]&selector_enabled,
r_1_addr[5]&r_0_addr[3]&selector_enabled,
r_1_addr[5]&r_0_addr[2]&selector_enabled,
r_1_addr[5]&r_0_addr[1]&selector_enabled,
r_1_addr[5]&r_0_addr[0]&selector_enabled,
r_1_addr[4]&r_0_addr[7]&selector_enabled,
r_1_addr[4]&r_0_addr[6]&selector_enabled,
r_1_addr[4]&r_0_addr[5]&selector_enabled,
r_1_addr[4]&r_0_addr[4]&selector_enabled,
r_1_addr[4]&r_0_addr[3]&selector_enabled,
r_1_addr[4]&r_0_addr[2]&selector_enabled,
r_1_addr[4]&r_0_addr[1]&selector_enabled,
r_1_addr[4]&r_0_addr[0]&selector_enabled,
r_1_addr[3]&r_0_addr[7]&selector_enabled,
r_1_addr[3]&r_0_addr[6]&selector_enabled,
r_1_addr[3]&r_0_addr[5]&selector_enabled,
r_1_addr[3]&r_0_addr[4]&selector_enabled,
r_1_addr[3]&r_0_addr[3]&selector_enabled,
r_1_addr[3]&r_0_addr[2]&selector_enabled,
r_1_addr[3]&r_0_addr[1]&selector_enabled,
r_1_addr[3]&r_0_addr[0]&selector_enabled,
r_1_addr[2]&r_0_addr[7]&selector_enabled,
r_1_addr[2]&r_0_addr[6]&selector_enabled,
r_1_addr[2]&r_0_addr[5]&selector_enabled,
r_1_addr[2]&r_0_addr[4]&selector_enabled,
r_1_addr[2]&r_0_addr[3]&selector_enabled,
r_1_addr[2]&r_0_addr[2]&selector_enabled,
r_1_addr[2]&r_0_addr[1]&selector_enabled,
r_1_addr[2]&r_0_addr[0]&selector_enabled,
r_1_addr[1]&r_0_addr[7]&selector_enabled,
r_1_addr[1]&r_0_addr[6]&selector_enabled,
r_1_addr[1]&r_0_addr[5]&selector_enabled,
r_1_addr[1]&r_0_addr[4]&selector_enabled,
r_1_addr[1]&r_0_addr[3]&selector_enabled,
r_1_addr[1]&r_0_addr[2]&selector_enabled,
r_1_addr[1]&r_0_addr[1]&selector_enabled,
r_1_addr[1]&r_0_addr[0]&selector_enabled,
r_1_addr[0]&r_0_addr[7]&selector_enabled,
r_1_addr[0]&r_0_addr[6]&selector_enabled,
r_1_addr[0]&r_0_addr[5]&selector_enabled,
r_1_addr[0]&r_0_addr[4]&selector_enabled,
r_1_addr[0]&r_0_addr[3]&selector_enabled,
r_1_addr[0]&r_0_addr[2]&selector_enabled,
r_1_addr[0]&r_0_addr[1]&selector_enabled,
r_1_addr[0]&r_0_addr[0]&selector_enabled};


endmodule
module memory_6

(input wire clk,
input wire write_en,
input wire[63:0] addr_selector_1,
input wire[63:0] addr_selector_2,
input wire[15:0] data_in,
output reg[15:0] data_out

);
reg[15:0] r_0_0;
reg[15:0] r_0_1;
reg[15:0] r_0_2;
reg[15:0] r_0_3;
reg[15:0] r_0_4;
reg[15:0] r_0_5;
reg[15:0] r_0_6;
reg[15:0] r_0_7;
reg[15:0] r_0_8;
reg[15:0] r_0_9;
reg[15:0] r_0_10;
reg[15:0] r_0_11;
reg[15:0] r_0_12;
reg[15:0] r_0_13;
reg[15:0] r_0_14;
reg[15:0] r_0_15;
reg[15:0] r_0_16;
reg[15:0] r_0_17;
reg[15:0] r_0_18;
reg[15:0] r_0_19;
reg[15:0] r_0_20;
reg[15:0] r_0_21;
reg[15:0] r_0_22;
reg[15:0] r_0_23;
reg[15:0] r_0_24;
reg[15:0] r_0_25;
reg[15:0] r_0_26;
reg[15:0] r_0_27;
reg[15:0] r_0_28;
reg[15:0] r_0_29;
reg[15:0] r_0_30;
reg[15:0] r_0_31;
reg[15:0] r_0_32;
reg[15:0] r_0_33;
reg[15:0] r_0_34;
reg[15:0] r_0_35;
reg[15:0] r_0_36;
reg[15:0] r_0_37;
reg[15:0] r_0_38;
reg[15:0] r_0_39;
reg[15:0] r_0_40;
reg[15:0] r_0_41;
reg[15:0] r_0_42;
reg[15:0] r_0_43;
reg[15:0] r_0_44;
reg[15:0] r_0_45;
reg[15:0] r_0_46;
reg[15:0] r_0_47;
reg[15:0] r_0_48;
reg[15:0] r_0_49;
reg[15:0] r_0_50;
reg[15:0] r_0_51;
reg[15:0] r_0_52;
reg[15:0] r_0_53;
reg[15:0] r_0_54;
reg[15:0] r_0_55;
reg[15:0] r_0_56;
reg[15:0] r_0_57;
reg[15:0] r_0_58;
reg[15:0] r_0_59;
reg[15:0] r_0_60;
reg[15:0] r_0_61;
reg[15:0] r_0_62;
reg[15:0] r_0_63;
reg[15:0] r_1_0;
reg[15:0] r_1_1;
reg[15:0] r_1_2;
reg[15:0] r_1_3;
reg[15:0] r_1_4;
reg[15:0] r_1_5;
reg[15:0] r_1_6;
reg[15:0] r_1_7;
reg[15:0] r_1_8;
reg[15:0] r_1_9;
reg[15:0] r_1_10;
reg[15:0] r_1_11;
reg[15:0] r_1_12;
reg[15:0] r_1_13;
reg[15:0] r_1_14;
reg[15:0] r_1_15;
reg[15:0] r_1_16;
reg[15:0] r_1_17;
reg[15:0] r_1_18;
reg[15:0] r_1_19;
reg[15:0] r_1_20;
reg[15:0] r_1_21;
reg[15:0] r_1_22;
reg[15:0] r_1_23;
reg[15:0] r_1_24;
reg[15:0] r_1_25;
reg[15:0] r_1_26;
reg[15:0] r_1_27;
reg[15:0] r_1_28;
reg[15:0] r_1_29;
reg[15:0] r_1_30;
reg[15:0] r_1_31;
reg[15:0] r_1_32;
reg[15:0] r_1_33;
reg[15:0] r_1_34;
reg[15:0] r_1_35;
reg[15:0] r_1_36;
reg[15:0] r_1_37;
reg[15:0] r_1_38;
reg[15:0] r_1_39;
reg[15:0] r_1_40;
reg[15:0] r_1_41;
reg[15:0] r_1_42;
reg[15:0] r_1_43;
reg[15:0] r_1_44;
reg[15:0] r_1_45;
reg[15:0] r_1_46;
reg[15:0] r_1_47;
reg[15:0] r_1_48;
reg[15:0] r_1_49;
reg[15:0] r_1_50;
reg[15:0] r_1_51;
reg[15:0] r_1_52;
reg[15:0] r_1_53;
reg[15:0] r_1_54;
reg[15:0] r_1_55;
reg[15:0] r_1_56;
reg[15:0] r_1_57;
reg[15:0] r_1_58;
reg[15:0] r_1_59;
reg[15:0] r_1_60;
reg[15:0] r_1_61;
reg[15:0] r_1_62;
reg[15:0] r_1_63;
reg[15:0] r_2_0;
reg[15:0] r_2_1;
reg[15:0] r_2_2;
reg[15:0] r_2_3;
reg[15:0] r_2_4;
reg[15:0] r_2_5;
reg[15:0] r_2_6;
reg[15:0] r_2_7;
reg[15:0] r_2_8;
reg[15:0] r_2_9;
reg[15:0] r_2_10;
reg[15:0] r_2_11;
reg[15:0] r_2_12;
reg[15:0] r_2_13;
reg[15:0] r_2_14;
reg[15:0] r_2_15;
reg[15:0] r_2_16;
reg[15:0] r_2_17;
reg[15:0] r_2_18;
reg[15:0] r_2_19;
reg[15:0] r_2_20;
reg[15:0] r_2_21;
reg[15:0] r_2_22;
reg[15:0] r_2_23;
reg[15:0] r_2_24;
reg[15:0] r_2_25;
reg[15:0] r_2_26;
reg[15:0] r_2_27;
reg[15:0] r_2_28;
reg[15:0] r_2_29;
reg[15:0] r_2_30;
reg[15:0] r_2_31;
reg[15:0] r_2_32;
reg[15:0] r_2_33;
reg[15:0] r_2_34;
reg[15:0] r_2_35;
reg[15:0] r_2_36;
reg[15:0] r_2_37;
reg[15:0] r_2_38;
reg[15:0] r_2_39;
reg[15:0] r_2_40;
reg[15:0] r_2_41;
reg[15:0] r_2_42;
reg[15:0] r_2_43;
reg[15:0] r_2_44;
reg[15:0] r_2_45;
reg[15:0] r_2_46;
reg[15:0] r_2_47;
reg[15:0] r_2_48;
reg[15:0] r_2_49;
reg[15:0] r_2_50;
reg[15:0] r_2_51;
reg[15:0] r_2_52;
reg[15:0] r_2_53;
reg[15:0] r_2_54;
reg[15:0] r_2_55;
reg[15:0] r_2_56;
reg[15:0] r_2_57;
reg[15:0] r_2_58;
reg[15:0] r_2_59;
reg[15:0] r_2_60;
reg[15:0] r_2_61;
reg[15:0] r_2_62;
reg[15:0] r_2_63;
reg[15:0] r_3_0;
reg[15:0] r_3_1;
reg[15:0] r_3_2;
reg[15:0] r_3_3;
reg[15:0] r_3_4;
reg[15:0] r_3_5;
reg[15:0] r_3_6;
reg[15:0] r_3_7;
reg[15:0] r_3_8;
reg[15:0] r_3_9;
reg[15:0] r_3_10;
reg[15:0] r_3_11;
reg[15:0] r_3_12;
reg[15:0] r_3_13;
reg[15:0] r_3_14;
reg[15:0] r_3_15;
reg[15:0] r_3_16;
reg[15:0] r_3_17;
reg[15:0] r_3_18;
reg[15:0] r_3_19;
reg[15:0] r_3_20;
reg[15:0] r_3_21;
reg[15:0] r_3_22;
reg[15:0] r_3_23;
reg[15:0] r_3_24;
reg[15:0] r_3_25;
reg[15:0] r_3_26;
reg[15:0] r_3_27;
reg[15:0] r_3_28;
reg[15:0] r_3_29;
reg[15:0] r_3_30;
reg[15:0] r_3_31;
reg[15:0] r_3_32;
reg[15:0] r_3_33;
reg[15:0] r_3_34;
reg[15:0] r_3_35;
reg[15:0] r_3_36;
reg[15:0] r_3_37;
reg[15:0] r_3_38;
reg[15:0] r_3_39;
reg[15:0] r_3_40;
reg[15:0] r_3_41;
reg[15:0] r_3_42;
reg[15:0] r_3_43;
reg[15:0] r_3_44;
reg[15:0] r_3_45;
reg[15:0] r_3_46;
reg[15:0] r_3_47;
reg[15:0] r_3_48;
reg[15:0] r_3_49;
reg[15:0] r_3_50;
reg[15:0] r_3_51;
reg[15:0] r_3_52;
reg[15:0] r_3_53;
reg[15:0] r_3_54;
reg[15:0] r_3_55;
reg[15:0] r_3_56;
reg[15:0] r_3_57;
reg[15:0] r_3_58;
reg[15:0] r_3_59;
reg[15:0] r_3_60;
reg[15:0] r_3_61;
reg[15:0] r_3_62;
reg[15:0] r_3_63;
reg[15:0] r_4_0;
reg[15:0] r_4_1;
reg[15:0] r_4_2;
reg[15:0] r_4_3;
reg[15:0] r_4_4;
reg[15:0] r_4_5;
reg[15:0] r_4_6;
reg[15:0] r_4_7;
reg[15:0] r_4_8;
reg[15:0] r_4_9;
reg[15:0] r_4_10;
reg[15:0] r_4_11;
reg[15:0] r_4_12;
reg[15:0] r_4_13;
reg[15:0] r_4_14;
reg[15:0] r_4_15;
reg[15:0] r_4_16;
reg[15:0] r_4_17;
reg[15:0] r_4_18;
reg[15:0] r_4_19;
reg[15:0] r_4_20;
reg[15:0] r_4_21;
reg[15:0] r_4_22;
reg[15:0] r_4_23;
reg[15:0] r_4_24;
reg[15:0] r_4_25;
reg[15:0] r_4_26;
reg[15:0] r_4_27;
reg[15:0] r_4_28;
reg[15:0] r_4_29;
reg[15:0] r_4_30;
reg[15:0] r_4_31;
reg[15:0] r_4_32;
reg[15:0] r_4_33;
reg[15:0] r_4_34;
reg[15:0] r_4_35;
reg[15:0] r_4_36;
reg[15:0] r_4_37;
reg[15:0] r_4_38;
reg[15:0] r_4_39;
reg[15:0] r_4_40;
reg[15:0] r_4_41;
reg[15:0] r_4_42;
reg[15:0] r_4_43;
reg[15:0] r_4_44;
reg[15:0] r_4_45;
reg[15:0] r_4_46;
reg[15:0] r_4_47;
reg[15:0] r_4_48;
reg[15:0] r_4_49;
reg[15:0] r_4_50;
reg[15:0] r_4_51;
reg[15:0] r_4_52;
reg[15:0] r_4_53;
reg[15:0] r_4_54;
reg[15:0] r_4_55;
reg[15:0] r_4_56;
reg[15:0] r_4_57;
reg[15:0] r_4_58;
reg[15:0] r_4_59;
reg[15:0] r_4_60;
reg[15:0] r_4_61;
reg[15:0] r_4_62;
reg[15:0] r_4_63;
reg[15:0] r_5_0;
reg[15:0] r_5_1;
reg[15:0] r_5_2;
reg[15:0] r_5_3;
reg[15:0] r_5_4;
reg[15:0] r_5_5;
reg[15:0] r_5_6;
reg[15:0] r_5_7;
reg[15:0] r_5_8;
reg[15:0] r_5_9;
reg[15:0] r_5_10;
reg[15:0] r_5_11;
reg[15:0] r_5_12;
reg[15:0] r_5_13;
reg[15:0] r_5_14;
reg[15:0] r_5_15;
reg[15:0] r_5_16;
reg[15:0] r_5_17;
reg[15:0] r_5_18;
reg[15:0] r_5_19;
reg[15:0] r_5_20;
reg[15:0] r_5_21;
reg[15:0] r_5_22;
reg[15:0] r_5_23;
reg[15:0] r_5_24;
reg[15:0] r_5_25;
reg[15:0] r_5_26;
reg[15:0] r_5_27;
reg[15:0] r_5_28;
reg[15:0] r_5_29;
reg[15:0] r_5_30;
reg[15:0] r_5_31;
reg[15:0] r_5_32;
reg[15:0] r_5_33;
reg[15:0] r_5_34;
reg[15:0] r_5_35;
reg[15:0] r_5_36;
reg[15:0] r_5_37;
reg[15:0] r_5_38;
reg[15:0] r_5_39;
reg[15:0] r_5_40;
reg[15:0] r_5_41;
reg[15:0] r_5_42;
reg[15:0] r_5_43;
reg[15:0] r_5_44;
reg[15:0] r_5_45;
reg[15:0] r_5_46;
reg[15:0] r_5_47;
reg[15:0] r_5_48;
reg[15:0] r_5_49;
reg[15:0] r_5_50;
reg[15:0] r_5_51;
reg[15:0] r_5_52;
reg[15:0] r_5_53;
reg[15:0] r_5_54;
reg[15:0] r_5_55;
reg[15:0] r_5_56;
reg[15:0] r_5_57;
reg[15:0] r_5_58;
reg[15:0] r_5_59;
reg[15:0] r_5_60;
reg[15:0] r_5_61;
reg[15:0] r_5_62;
reg[15:0] r_5_63;
reg[15:0] r_6_0;
reg[15:0] r_6_1;
reg[15:0] r_6_2;
reg[15:0] r_6_3;
reg[15:0] r_6_4;
reg[15:0] r_6_5;
reg[15:0] r_6_6;
reg[15:0] r_6_7;
reg[15:0] r_6_8;
reg[15:0] r_6_9;
reg[15:0] r_6_10;
reg[15:0] r_6_11;
reg[15:0] r_6_12;
reg[15:0] r_6_13;
reg[15:0] r_6_14;
reg[15:0] r_6_15;
reg[15:0] r_6_16;
reg[15:0] r_6_17;
reg[15:0] r_6_18;
reg[15:0] r_6_19;
reg[15:0] r_6_20;
reg[15:0] r_6_21;
reg[15:0] r_6_22;
reg[15:0] r_6_23;
reg[15:0] r_6_24;
reg[15:0] r_6_25;
reg[15:0] r_6_26;
reg[15:0] r_6_27;
reg[15:0] r_6_28;
reg[15:0] r_6_29;
reg[15:0] r_6_30;
reg[15:0] r_6_31;
reg[15:0] r_6_32;
reg[15:0] r_6_33;
reg[15:0] r_6_34;
reg[15:0] r_6_35;
reg[15:0] r_6_36;
reg[15:0] r_6_37;
reg[15:0] r_6_38;
reg[15:0] r_6_39;
reg[15:0] r_6_40;
reg[15:0] r_6_41;
reg[15:0] r_6_42;
reg[15:0] r_6_43;
reg[15:0] r_6_44;
reg[15:0] r_6_45;
reg[15:0] r_6_46;
reg[15:0] r_6_47;
reg[15:0] r_6_48;
reg[15:0] r_6_49;
reg[15:0] r_6_50;
reg[15:0] r_6_51;
reg[15:0] r_6_52;
reg[15:0] r_6_53;
reg[15:0] r_6_54;
reg[15:0] r_6_55;
reg[15:0] r_6_56;
reg[15:0] r_6_57;
reg[15:0] r_6_58;
reg[15:0] r_6_59;
reg[15:0] r_6_60;
reg[15:0] r_6_61;
reg[15:0] r_6_62;
reg[15:0] r_6_63;
reg[15:0] r_7_0;
reg[15:0] r_7_1;
reg[15:0] r_7_2;
reg[15:0] r_7_3;
reg[15:0] r_7_4;
reg[15:0] r_7_5;
reg[15:0] r_7_6;
reg[15:0] r_7_7;
reg[15:0] r_7_8;
reg[15:0] r_7_9;
reg[15:0] r_7_10;
reg[15:0] r_7_11;
reg[15:0] r_7_12;
reg[15:0] r_7_13;
reg[15:0] r_7_14;
reg[15:0] r_7_15;
reg[15:0] r_7_16;
reg[15:0] r_7_17;
reg[15:0] r_7_18;
reg[15:0] r_7_19;
reg[15:0] r_7_20;
reg[15:0] r_7_21;
reg[15:0] r_7_22;
reg[15:0] r_7_23;
reg[15:0] r_7_24;
reg[15:0] r_7_25;
reg[15:0] r_7_26;
reg[15:0] r_7_27;
reg[15:0] r_7_28;
reg[15:0] r_7_29;
reg[15:0] r_7_30;
reg[15:0] r_7_31;
reg[15:0] r_7_32;
reg[15:0] r_7_33;
reg[15:0] r_7_34;
reg[15:0] r_7_35;
reg[15:0] r_7_36;
reg[15:0] r_7_37;
reg[15:0] r_7_38;
reg[15:0] r_7_39;
reg[15:0] r_7_40;
reg[15:0] r_7_41;
reg[15:0] r_7_42;
reg[15:0] r_7_43;
reg[15:0] r_7_44;
reg[15:0] r_7_45;
reg[15:0] r_7_46;
reg[15:0] r_7_47;
reg[15:0] r_7_48;
reg[15:0] r_7_49;
reg[15:0] r_7_50;
reg[15:0] r_7_51;
reg[15:0] r_7_52;
reg[15:0] r_7_53;
reg[15:0] r_7_54;
reg[15:0] r_7_55;
reg[15:0] r_7_56;
reg[15:0] r_7_57;
reg[15:0] r_7_58;
reg[15:0] r_7_59;
reg[15:0] r_7_60;
reg[15:0] r_7_61;
reg[15:0] r_7_62;
reg[15:0] r_7_63;
reg[15:0] r_8_0;
reg[15:0] r_8_1;
reg[15:0] r_8_2;
reg[15:0] r_8_3;
reg[15:0] r_8_4;
reg[15:0] r_8_5;
reg[15:0] r_8_6;
reg[15:0] r_8_7;
reg[15:0] r_8_8;
reg[15:0] r_8_9;
reg[15:0] r_8_10;
reg[15:0] r_8_11;
reg[15:0] r_8_12;
reg[15:0] r_8_13;
reg[15:0] r_8_14;
reg[15:0] r_8_15;
reg[15:0] r_8_16;
reg[15:0] r_8_17;
reg[15:0] r_8_18;
reg[15:0] r_8_19;
reg[15:0] r_8_20;
reg[15:0] r_8_21;
reg[15:0] r_8_22;
reg[15:0] r_8_23;
reg[15:0] r_8_24;
reg[15:0] r_8_25;
reg[15:0] r_8_26;
reg[15:0] r_8_27;
reg[15:0] r_8_28;
reg[15:0] r_8_29;
reg[15:0] r_8_30;
reg[15:0] r_8_31;
reg[15:0] r_8_32;
reg[15:0] r_8_33;
reg[15:0] r_8_34;
reg[15:0] r_8_35;
reg[15:0] r_8_36;
reg[15:0] r_8_37;
reg[15:0] r_8_38;
reg[15:0] r_8_39;
reg[15:0] r_8_40;
reg[15:0] r_8_41;
reg[15:0] r_8_42;
reg[15:0] r_8_43;
reg[15:0] r_8_44;
reg[15:0] r_8_45;
reg[15:0] r_8_46;
reg[15:0] r_8_47;
reg[15:0] r_8_48;
reg[15:0] r_8_49;
reg[15:0] r_8_50;
reg[15:0] r_8_51;
reg[15:0] r_8_52;
reg[15:0] r_8_53;
reg[15:0] r_8_54;
reg[15:0] r_8_55;
reg[15:0] r_8_56;
reg[15:0] r_8_57;
reg[15:0] r_8_58;
reg[15:0] r_8_59;
reg[15:0] r_8_60;
reg[15:0] r_8_61;
reg[15:0] r_8_62;
reg[15:0] r_8_63;
reg[15:0] r_9_0;
reg[15:0] r_9_1;
reg[15:0] r_9_2;
reg[15:0] r_9_3;
reg[15:0] r_9_4;
reg[15:0] r_9_5;
reg[15:0] r_9_6;
reg[15:0] r_9_7;
reg[15:0] r_9_8;
reg[15:0] r_9_9;
reg[15:0] r_9_10;
reg[15:0] r_9_11;
reg[15:0] r_9_12;
reg[15:0] r_9_13;
reg[15:0] r_9_14;
reg[15:0] r_9_15;
reg[15:0] r_9_16;
reg[15:0] r_9_17;
reg[15:0] r_9_18;
reg[15:0] r_9_19;
reg[15:0] r_9_20;
reg[15:0] r_9_21;
reg[15:0] r_9_22;
reg[15:0] r_9_23;
reg[15:0] r_9_24;
reg[15:0] r_9_25;
reg[15:0] r_9_26;
reg[15:0] r_9_27;
reg[15:0] r_9_28;
reg[15:0] r_9_29;
reg[15:0] r_9_30;
reg[15:0] r_9_31;
reg[15:0] r_9_32;
reg[15:0] r_9_33;
reg[15:0] r_9_34;
reg[15:0] r_9_35;
reg[15:0] r_9_36;
reg[15:0] r_9_37;
reg[15:0] r_9_38;
reg[15:0] r_9_39;
reg[15:0] r_9_40;
reg[15:0] r_9_41;
reg[15:0] r_9_42;
reg[15:0] r_9_43;
reg[15:0] r_9_44;
reg[15:0] r_9_45;
reg[15:0] r_9_46;
reg[15:0] r_9_47;
reg[15:0] r_9_48;
reg[15:0] r_9_49;
reg[15:0] r_9_50;
reg[15:0] r_9_51;
reg[15:0] r_9_52;
reg[15:0] r_9_53;
reg[15:0] r_9_54;
reg[15:0] r_9_55;
reg[15:0] r_9_56;
reg[15:0] r_9_57;
reg[15:0] r_9_58;
reg[15:0] r_9_59;
reg[15:0] r_9_60;
reg[15:0] r_9_61;
reg[15:0] r_9_62;
reg[15:0] r_9_63;
reg[15:0] r_10_0;
reg[15:0] r_10_1;
reg[15:0] r_10_2;
reg[15:0] r_10_3;
reg[15:0] r_10_4;
reg[15:0] r_10_5;
reg[15:0] r_10_6;
reg[15:0] r_10_7;
reg[15:0] r_10_8;
reg[15:0] r_10_9;
reg[15:0] r_10_10;
reg[15:0] r_10_11;
reg[15:0] r_10_12;
reg[15:0] r_10_13;
reg[15:0] r_10_14;
reg[15:0] r_10_15;
reg[15:0] r_10_16;
reg[15:0] r_10_17;
reg[15:0] r_10_18;
reg[15:0] r_10_19;
reg[15:0] r_10_20;
reg[15:0] r_10_21;
reg[15:0] r_10_22;
reg[15:0] r_10_23;
reg[15:0] r_10_24;
reg[15:0] r_10_25;
reg[15:0] r_10_26;
reg[15:0] r_10_27;
reg[15:0] r_10_28;
reg[15:0] r_10_29;
reg[15:0] r_10_30;
reg[15:0] r_10_31;
reg[15:0] r_10_32;
reg[15:0] r_10_33;
reg[15:0] r_10_34;
reg[15:0] r_10_35;
reg[15:0] r_10_36;
reg[15:0] r_10_37;
reg[15:0] r_10_38;
reg[15:0] r_10_39;
reg[15:0] r_10_40;
reg[15:0] r_10_41;
reg[15:0] r_10_42;
reg[15:0] r_10_43;
reg[15:0] r_10_44;
reg[15:0] r_10_45;
reg[15:0] r_10_46;
reg[15:0] r_10_47;
reg[15:0] r_10_48;
reg[15:0] r_10_49;
reg[15:0] r_10_50;
reg[15:0] r_10_51;
reg[15:0] r_10_52;
reg[15:0] r_10_53;
reg[15:0] r_10_54;
reg[15:0] r_10_55;
reg[15:0] r_10_56;
reg[15:0] r_10_57;
reg[15:0] r_10_58;
reg[15:0] r_10_59;
reg[15:0] r_10_60;
reg[15:0] r_10_61;
reg[15:0] r_10_62;
reg[15:0] r_10_63;
reg[15:0] r_11_0;
reg[15:0] r_11_1;
reg[15:0] r_11_2;
reg[15:0] r_11_3;
reg[15:0] r_11_4;
reg[15:0] r_11_5;
reg[15:0] r_11_6;
reg[15:0] r_11_7;
reg[15:0] r_11_8;
reg[15:0] r_11_9;
reg[15:0] r_11_10;
reg[15:0] r_11_11;
reg[15:0] r_11_12;
reg[15:0] r_11_13;
reg[15:0] r_11_14;
reg[15:0] r_11_15;
reg[15:0] r_11_16;
reg[15:0] r_11_17;
reg[15:0] r_11_18;
reg[15:0] r_11_19;
reg[15:0] r_11_20;
reg[15:0] r_11_21;
reg[15:0] r_11_22;
reg[15:0] r_11_23;
reg[15:0] r_11_24;
reg[15:0] r_11_25;
reg[15:0] r_11_26;
reg[15:0] r_11_27;
reg[15:0] r_11_28;
reg[15:0] r_11_29;
reg[15:0] r_11_30;
reg[15:0] r_11_31;
reg[15:0] r_11_32;
reg[15:0] r_11_33;
reg[15:0] r_11_34;
reg[15:0] r_11_35;
reg[15:0] r_11_36;
reg[15:0] r_11_37;
reg[15:0] r_11_38;
reg[15:0] r_11_39;
reg[15:0] r_11_40;
reg[15:0] r_11_41;
reg[15:0] r_11_42;
reg[15:0] r_11_43;
reg[15:0] r_11_44;
reg[15:0] r_11_45;
reg[15:0] r_11_46;
reg[15:0] r_11_47;
reg[15:0] r_11_48;
reg[15:0] r_11_49;
reg[15:0] r_11_50;
reg[15:0] r_11_51;
reg[15:0] r_11_52;
reg[15:0] r_11_53;
reg[15:0] r_11_54;
reg[15:0] r_11_55;
reg[15:0] r_11_56;
reg[15:0] r_11_57;
reg[15:0] r_11_58;
reg[15:0] r_11_59;
reg[15:0] r_11_60;
reg[15:0] r_11_61;
reg[15:0] r_11_62;
reg[15:0] r_11_63;
reg[15:0] r_12_0;
reg[15:0] r_12_1;
reg[15:0] r_12_2;
reg[15:0] r_12_3;
reg[15:0] r_12_4;
reg[15:0] r_12_5;
reg[15:0] r_12_6;
reg[15:0] r_12_7;
reg[15:0] r_12_8;
reg[15:0] r_12_9;
reg[15:0] r_12_10;
reg[15:0] r_12_11;
reg[15:0] r_12_12;
reg[15:0] r_12_13;
reg[15:0] r_12_14;
reg[15:0] r_12_15;
reg[15:0] r_12_16;
reg[15:0] r_12_17;
reg[15:0] r_12_18;
reg[15:0] r_12_19;
reg[15:0] r_12_20;
reg[15:0] r_12_21;
reg[15:0] r_12_22;
reg[15:0] r_12_23;
reg[15:0] r_12_24;
reg[15:0] r_12_25;
reg[15:0] r_12_26;
reg[15:0] r_12_27;
reg[15:0] r_12_28;
reg[15:0] r_12_29;
reg[15:0] r_12_30;
reg[15:0] r_12_31;
reg[15:0] r_12_32;
reg[15:0] r_12_33;
reg[15:0] r_12_34;
reg[15:0] r_12_35;
reg[15:0] r_12_36;
reg[15:0] r_12_37;
reg[15:0] r_12_38;
reg[15:0] r_12_39;
reg[15:0] r_12_40;
reg[15:0] r_12_41;
reg[15:0] r_12_42;
reg[15:0] r_12_43;
reg[15:0] r_12_44;
reg[15:0] r_12_45;
reg[15:0] r_12_46;
reg[15:0] r_12_47;
reg[15:0] r_12_48;
reg[15:0] r_12_49;
reg[15:0] r_12_50;
reg[15:0] r_12_51;
reg[15:0] r_12_52;
reg[15:0] r_12_53;
reg[15:0] r_12_54;
reg[15:0] r_12_55;
reg[15:0] r_12_56;
reg[15:0] r_12_57;
reg[15:0] r_12_58;
reg[15:0] r_12_59;
reg[15:0] r_12_60;
reg[15:0] r_12_61;
reg[15:0] r_12_62;
reg[15:0] r_12_63;
reg[15:0] r_13_0;
reg[15:0] r_13_1;
reg[15:0] r_13_2;
reg[15:0] r_13_3;
reg[15:0] r_13_4;
reg[15:0] r_13_5;
reg[15:0] r_13_6;
reg[15:0] r_13_7;
reg[15:0] r_13_8;
reg[15:0] r_13_9;
reg[15:0] r_13_10;
reg[15:0] r_13_11;
reg[15:0] r_13_12;
reg[15:0] r_13_13;
reg[15:0] r_13_14;
reg[15:0] r_13_15;
reg[15:0] r_13_16;
reg[15:0] r_13_17;
reg[15:0] r_13_18;
reg[15:0] r_13_19;
reg[15:0] r_13_20;
reg[15:0] r_13_21;
reg[15:0] r_13_22;
reg[15:0] r_13_23;
reg[15:0] r_13_24;
reg[15:0] r_13_25;
reg[15:0] r_13_26;
reg[15:0] r_13_27;
reg[15:0] r_13_28;
reg[15:0] r_13_29;
reg[15:0] r_13_30;
reg[15:0] r_13_31;
reg[15:0] r_13_32;
reg[15:0] r_13_33;
reg[15:0] r_13_34;
reg[15:0] r_13_35;
reg[15:0] r_13_36;
reg[15:0] r_13_37;
reg[15:0] r_13_38;
reg[15:0] r_13_39;
reg[15:0] r_13_40;
reg[15:0] r_13_41;
reg[15:0] r_13_42;
reg[15:0] r_13_43;
reg[15:0] r_13_44;
reg[15:0] r_13_45;
reg[15:0] r_13_46;
reg[15:0] r_13_47;
reg[15:0] r_13_48;
reg[15:0] r_13_49;
reg[15:0] r_13_50;
reg[15:0] r_13_51;
reg[15:0] r_13_52;
reg[15:0] r_13_53;
reg[15:0] r_13_54;
reg[15:0] r_13_55;
reg[15:0] r_13_56;
reg[15:0] r_13_57;
reg[15:0] r_13_58;
reg[15:0] r_13_59;
reg[15:0] r_13_60;
reg[15:0] r_13_61;
reg[15:0] r_13_62;
reg[15:0] r_13_63;
reg[15:0] r_14_0;
reg[15:0] r_14_1;
reg[15:0] r_14_2;
reg[15:0] r_14_3;
reg[15:0] r_14_4;
reg[15:0] r_14_5;
reg[15:0] r_14_6;
reg[15:0] r_14_7;
reg[15:0] r_14_8;
reg[15:0] r_14_9;
reg[15:0] r_14_10;
reg[15:0] r_14_11;
reg[15:0] r_14_12;
reg[15:0] r_14_13;
reg[15:0] r_14_14;
reg[15:0] r_14_15;
reg[15:0] r_14_16;
reg[15:0] r_14_17;
reg[15:0] r_14_18;
reg[15:0] r_14_19;
reg[15:0] r_14_20;
reg[15:0] r_14_21;
reg[15:0] r_14_22;
reg[15:0] r_14_23;
reg[15:0] r_14_24;
reg[15:0] r_14_25;
reg[15:0] r_14_26;
reg[15:0] r_14_27;
reg[15:0] r_14_28;
reg[15:0] r_14_29;
reg[15:0] r_14_30;
reg[15:0] r_14_31;
reg[15:0] r_14_32;
reg[15:0] r_14_33;
reg[15:0] r_14_34;
reg[15:0] r_14_35;
reg[15:0] r_14_36;
reg[15:0] r_14_37;
reg[15:0] r_14_38;
reg[15:0] r_14_39;
reg[15:0] r_14_40;
reg[15:0] r_14_41;
reg[15:0] r_14_42;
reg[15:0] r_14_43;
reg[15:0] r_14_44;
reg[15:0] r_14_45;
reg[15:0] r_14_46;
reg[15:0] r_14_47;
reg[15:0] r_14_48;
reg[15:0] r_14_49;
reg[15:0] r_14_50;
reg[15:0] r_14_51;
reg[15:0] r_14_52;
reg[15:0] r_14_53;
reg[15:0] r_14_54;
reg[15:0] r_14_55;
reg[15:0] r_14_56;
reg[15:0] r_14_57;
reg[15:0] r_14_58;
reg[15:0] r_14_59;
reg[15:0] r_14_60;
reg[15:0] r_14_61;
reg[15:0] r_14_62;
reg[15:0] r_14_63;
reg[15:0] r_15_0;
reg[15:0] r_15_1;
reg[15:0] r_15_2;
reg[15:0] r_15_3;
reg[15:0] r_15_4;
reg[15:0] r_15_5;
reg[15:0] r_15_6;
reg[15:0] r_15_7;
reg[15:0] r_15_8;
reg[15:0] r_15_9;
reg[15:0] r_15_10;
reg[15:0] r_15_11;
reg[15:0] r_15_12;
reg[15:0] r_15_13;
reg[15:0] r_15_14;
reg[15:0] r_15_15;
reg[15:0] r_15_16;
reg[15:0] r_15_17;
reg[15:0] r_15_18;
reg[15:0] r_15_19;
reg[15:0] r_15_20;
reg[15:0] r_15_21;
reg[15:0] r_15_22;
reg[15:0] r_15_23;
reg[15:0] r_15_24;
reg[15:0] r_15_25;
reg[15:0] r_15_26;
reg[15:0] r_15_27;
reg[15:0] r_15_28;
reg[15:0] r_15_29;
reg[15:0] r_15_30;
reg[15:0] r_15_31;
reg[15:0] r_15_32;
reg[15:0] r_15_33;
reg[15:0] r_15_34;
reg[15:0] r_15_35;
reg[15:0] r_15_36;
reg[15:0] r_15_37;
reg[15:0] r_15_38;
reg[15:0] r_15_39;
reg[15:0] r_15_40;
reg[15:0] r_15_41;
reg[15:0] r_15_42;
reg[15:0] r_15_43;
reg[15:0] r_15_44;
reg[15:0] r_15_45;
reg[15:0] r_15_46;
reg[15:0] r_15_47;
reg[15:0] r_15_48;
reg[15:0] r_15_49;
reg[15:0] r_15_50;
reg[15:0] r_15_51;
reg[15:0] r_15_52;
reg[15:0] r_15_53;
reg[15:0] r_15_54;
reg[15:0] r_15_55;
reg[15:0] r_15_56;
reg[15:0] r_15_57;
reg[15:0] r_15_58;
reg[15:0] r_15_59;
reg[15:0] r_15_60;
reg[15:0] r_15_61;
reg[15:0] r_15_62;
reg[15:0] r_15_63;
reg[15:0] r_16_0;
reg[15:0] r_16_1;
reg[15:0] r_16_2;
reg[15:0] r_16_3;
reg[15:0] r_16_4;
reg[15:0] r_16_5;
reg[15:0] r_16_6;
reg[15:0] r_16_7;
reg[15:0] r_16_8;
reg[15:0] r_16_9;
reg[15:0] r_16_10;
reg[15:0] r_16_11;
reg[15:0] r_16_12;
reg[15:0] r_16_13;
reg[15:0] r_16_14;
reg[15:0] r_16_15;
reg[15:0] r_16_16;
reg[15:0] r_16_17;
reg[15:0] r_16_18;
reg[15:0] r_16_19;
reg[15:0] r_16_20;
reg[15:0] r_16_21;
reg[15:0] r_16_22;
reg[15:0] r_16_23;
reg[15:0] r_16_24;
reg[15:0] r_16_25;
reg[15:0] r_16_26;
reg[15:0] r_16_27;
reg[15:0] r_16_28;
reg[15:0] r_16_29;
reg[15:0] r_16_30;
reg[15:0] r_16_31;
reg[15:0] r_16_32;
reg[15:0] r_16_33;
reg[15:0] r_16_34;
reg[15:0] r_16_35;
reg[15:0] r_16_36;
reg[15:0] r_16_37;
reg[15:0] r_16_38;
reg[15:0] r_16_39;
reg[15:0] r_16_40;
reg[15:0] r_16_41;
reg[15:0] r_16_42;
reg[15:0] r_16_43;
reg[15:0] r_16_44;
reg[15:0] r_16_45;
reg[15:0] r_16_46;
reg[15:0] r_16_47;
reg[15:0] r_16_48;
reg[15:0] r_16_49;
reg[15:0] r_16_50;
reg[15:0] r_16_51;
reg[15:0] r_16_52;
reg[15:0] r_16_53;
reg[15:0] r_16_54;
reg[15:0] r_16_55;
reg[15:0] r_16_56;
reg[15:0] r_16_57;
reg[15:0] r_16_58;
reg[15:0] r_16_59;
reg[15:0] r_16_60;
reg[15:0] r_16_61;
reg[15:0] r_16_62;
reg[15:0] r_16_63;
reg[15:0] r_17_0;
reg[15:0] r_17_1;
reg[15:0] r_17_2;
reg[15:0] r_17_3;
reg[15:0] r_17_4;
reg[15:0] r_17_5;
reg[15:0] r_17_6;
reg[15:0] r_17_7;
reg[15:0] r_17_8;
reg[15:0] r_17_9;
reg[15:0] r_17_10;
reg[15:0] r_17_11;
reg[15:0] r_17_12;
reg[15:0] r_17_13;
reg[15:0] r_17_14;
reg[15:0] r_17_15;
reg[15:0] r_17_16;
reg[15:0] r_17_17;
reg[15:0] r_17_18;
reg[15:0] r_17_19;
reg[15:0] r_17_20;
reg[15:0] r_17_21;
reg[15:0] r_17_22;
reg[15:0] r_17_23;
reg[15:0] r_17_24;
reg[15:0] r_17_25;
reg[15:0] r_17_26;
reg[15:0] r_17_27;
reg[15:0] r_17_28;
reg[15:0] r_17_29;
reg[15:0] r_17_30;
reg[15:0] r_17_31;
reg[15:0] r_17_32;
reg[15:0] r_17_33;
reg[15:0] r_17_34;
reg[15:0] r_17_35;
reg[15:0] r_17_36;
reg[15:0] r_17_37;
reg[15:0] r_17_38;
reg[15:0] r_17_39;
reg[15:0] r_17_40;
reg[15:0] r_17_41;
reg[15:0] r_17_42;
reg[15:0] r_17_43;
reg[15:0] r_17_44;
reg[15:0] r_17_45;
reg[15:0] r_17_46;
reg[15:0] r_17_47;
reg[15:0] r_17_48;
reg[15:0] r_17_49;
reg[15:0] r_17_50;
reg[15:0] r_17_51;
reg[15:0] r_17_52;
reg[15:0] r_17_53;
reg[15:0] r_17_54;
reg[15:0] r_17_55;
reg[15:0] r_17_56;
reg[15:0] r_17_57;
reg[15:0] r_17_58;
reg[15:0] r_17_59;
reg[15:0] r_17_60;
reg[15:0] r_17_61;
reg[15:0] r_17_62;
reg[15:0] r_17_63;
reg[15:0] r_18_0;
reg[15:0] r_18_1;
reg[15:0] r_18_2;
reg[15:0] r_18_3;
reg[15:0] r_18_4;
reg[15:0] r_18_5;
reg[15:0] r_18_6;
reg[15:0] r_18_7;
reg[15:0] r_18_8;
reg[15:0] r_18_9;
reg[15:0] r_18_10;
reg[15:0] r_18_11;
reg[15:0] r_18_12;
reg[15:0] r_18_13;
reg[15:0] r_18_14;
reg[15:0] r_18_15;
reg[15:0] r_18_16;
reg[15:0] r_18_17;
reg[15:0] r_18_18;
reg[15:0] r_18_19;
reg[15:0] r_18_20;
reg[15:0] r_18_21;
reg[15:0] r_18_22;
reg[15:0] r_18_23;
reg[15:0] r_18_24;
reg[15:0] r_18_25;
reg[15:0] r_18_26;
reg[15:0] r_18_27;
reg[15:0] r_18_28;
reg[15:0] r_18_29;
reg[15:0] r_18_30;
reg[15:0] r_18_31;
reg[15:0] r_18_32;
reg[15:0] r_18_33;
reg[15:0] r_18_34;
reg[15:0] r_18_35;
reg[15:0] r_18_36;
reg[15:0] r_18_37;
reg[15:0] r_18_38;
reg[15:0] r_18_39;
reg[15:0] r_18_40;
reg[15:0] r_18_41;
reg[15:0] r_18_42;
reg[15:0] r_18_43;
reg[15:0] r_18_44;
reg[15:0] r_18_45;
reg[15:0] r_18_46;
reg[15:0] r_18_47;
reg[15:0] r_18_48;
reg[15:0] r_18_49;
reg[15:0] r_18_50;
reg[15:0] r_18_51;
reg[15:0] r_18_52;
reg[15:0] r_18_53;
reg[15:0] r_18_54;
reg[15:0] r_18_55;
reg[15:0] r_18_56;
reg[15:0] r_18_57;
reg[15:0] r_18_58;
reg[15:0] r_18_59;
reg[15:0] r_18_60;
reg[15:0] r_18_61;
reg[15:0] r_18_62;
reg[15:0] r_18_63;
reg[15:0] r_19_0;
reg[15:0] r_19_1;
reg[15:0] r_19_2;
reg[15:0] r_19_3;
reg[15:0] r_19_4;
reg[15:0] r_19_5;
reg[15:0] r_19_6;
reg[15:0] r_19_7;
reg[15:0] r_19_8;
reg[15:0] r_19_9;
reg[15:0] r_19_10;
reg[15:0] r_19_11;
reg[15:0] r_19_12;
reg[15:0] r_19_13;
reg[15:0] r_19_14;
reg[15:0] r_19_15;
reg[15:0] r_19_16;
reg[15:0] r_19_17;
reg[15:0] r_19_18;
reg[15:0] r_19_19;
reg[15:0] r_19_20;
reg[15:0] r_19_21;
reg[15:0] r_19_22;
reg[15:0] r_19_23;
reg[15:0] r_19_24;
reg[15:0] r_19_25;
reg[15:0] r_19_26;
reg[15:0] r_19_27;
reg[15:0] r_19_28;
reg[15:0] r_19_29;
reg[15:0] r_19_30;
reg[15:0] r_19_31;
reg[15:0] r_19_32;
reg[15:0] r_19_33;
reg[15:0] r_19_34;
reg[15:0] r_19_35;
reg[15:0] r_19_36;
reg[15:0] r_19_37;
reg[15:0] r_19_38;
reg[15:0] r_19_39;
reg[15:0] r_19_40;
reg[15:0] r_19_41;
reg[15:0] r_19_42;
reg[15:0] r_19_43;
reg[15:0] r_19_44;
reg[15:0] r_19_45;
reg[15:0] r_19_46;
reg[15:0] r_19_47;
reg[15:0] r_19_48;
reg[15:0] r_19_49;
reg[15:0] r_19_50;
reg[15:0] r_19_51;
reg[15:0] r_19_52;
reg[15:0] r_19_53;
reg[15:0] r_19_54;
reg[15:0] r_19_55;
reg[15:0] r_19_56;
reg[15:0] r_19_57;
reg[15:0] r_19_58;
reg[15:0] r_19_59;
reg[15:0] r_19_60;
reg[15:0] r_19_61;
reg[15:0] r_19_62;
reg[15:0] r_19_63;
reg[15:0] r_20_0;
reg[15:0] r_20_1;
reg[15:0] r_20_2;
reg[15:0] r_20_3;
reg[15:0] r_20_4;
reg[15:0] r_20_5;
reg[15:0] r_20_6;
reg[15:0] r_20_7;
reg[15:0] r_20_8;
reg[15:0] r_20_9;
reg[15:0] r_20_10;
reg[15:0] r_20_11;
reg[15:0] r_20_12;
reg[15:0] r_20_13;
reg[15:0] r_20_14;
reg[15:0] r_20_15;
reg[15:0] r_20_16;
reg[15:0] r_20_17;
reg[15:0] r_20_18;
reg[15:0] r_20_19;
reg[15:0] r_20_20;
reg[15:0] r_20_21;
reg[15:0] r_20_22;
reg[15:0] r_20_23;
reg[15:0] r_20_24;
reg[15:0] r_20_25;
reg[15:0] r_20_26;
reg[15:0] r_20_27;
reg[15:0] r_20_28;
reg[15:0] r_20_29;
reg[15:0] r_20_30;
reg[15:0] r_20_31;
reg[15:0] r_20_32;
reg[15:0] r_20_33;
reg[15:0] r_20_34;
reg[15:0] r_20_35;
reg[15:0] r_20_36;
reg[15:0] r_20_37;
reg[15:0] r_20_38;
reg[15:0] r_20_39;
reg[15:0] r_20_40;
reg[15:0] r_20_41;
reg[15:0] r_20_42;
reg[15:0] r_20_43;
reg[15:0] r_20_44;
reg[15:0] r_20_45;
reg[15:0] r_20_46;
reg[15:0] r_20_47;
reg[15:0] r_20_48;
reg[15:0] r_20_49;
reg[15:0] r_20_50;
reg[15:0] r_20_51;
reg[15:0] r_20_52;
reg[15:0] r_20_53;
reg[15:0] r_20_54;
reg[15:0] r_20_55;
reg[15:0] r_20_56;
reg[15:0] r_20_57;
reg[15:0] r_20_58;
reg[15:0] r_20_59;
reg[15:0] r_20_60;
reg[15:0] r_20_61;
reg[15:0] r_20_62;
reg[15:0] r_20_63;
reg[15:0] r_21_0;
reg[15:0] r_21_1;
reg[15:0] r_21_2;
reg[15:0] r_21_3;
reg[15:0] r_21_4;
reg[15:0] r_21_5;
reg[15:0] r_21_6;
reg[15:0] r_21_7;
reg[15:0] r_21_8;
reg[15:0] r_21_9;
reg[15:0] r_21_10;
reg[15:0] r_21_11;
reg[15:0] r_21_12;
reg[15:0] r_21_13;
reg[15:0] r_21_14;
reg[15:0] r_21_15;
reg[15:0] r_21_16;
reg[15:0] r_21_17;
reg[15:0] r_21_18;
reg[15:0] r_21_19;
reg[15:0] r_21_20;
reg[15:0] r_21_21;
reg[15:0] r_21_22;
reg[15:0] r_21_23;
reg[15:0] r_21_24;
reg[15:0] r_21_25;
reg[15:0] r_21_26;
reg[15:0] r_21_27;
reg[15:0] r_21_28;
reg[15:0] r_21_29;
reg[15:0] r_21_30;
reg[15:0] r_21_31;
reg[15:0] r_21_32;
reg[15:0] r_21_33;
reg[15:0] r_21_34;
reg[15:0] r_21_35;
reg[15:0] r_21_36;
reg[15:0] r_21_37;
reg[15:0] r_21_38;
reg[15:0] r_21_39;
reg[15:0] r_21_40;
reg[15:0] r_21_41;
reg[15:0] r_21_42;
reg[15:0] r_21_43;
reg[15:0] r_21_44;
reg[15:0] r_21_45;
reg[15:0] r_21_46;
reg[15:0] r_21_47;
reg[15:0] r_21_48;
reg[15:0] r_21_49;
reg[15:0] r_21_50;
reg[15:0] r_21_51;
reg[15:0] r_21_52;
reg[15:0] r_21_53;
reg[15:0] r_21_54;
reg[15:0] r_21_55;
reg[15:0] r_21_56;
reg[15:0] r_21_57;
reg[15:0] r_21_58;
reg[15:0] r_21_59;
reg[15:0] r_21_60;
reg[15:0] r_21_61;
reg[15:0] r_21_62;
reg[15:0] r_21_63;
reg[15:0] r_22_0;
reg[15:0] r_22_1;
reg[15:0] r_22_2;
reg[15:0] r_22_3;
reg[15:0] r_22_4;
reg[15:0] r_22_5;
reg[15:0] r_22_6;
reg[15:0] r_22_7;
reg[15:0] r_22_8;
reg[15:0] r_22_9;
reg[15:0] r_22_10;
reg[15:0] r_22_11;
reg[15:0] r_22_12;
reg[15:0] r_22_13;
reg[15:0] r_22_14;
reg[15:0] r_22_15;
reg[15:0] r_22_16;
reg[15:0] r_22_17;
reg[15:0] r_22_18;
reg[15:0] r_22_19;
reg[15:0] r_22_20;
reg[15:0] r_22_21;
reg[15:0] r_22_22;
reg[15:0] r_22_23;
reg[15:0] r_22_24;
reg[15:0] r_22_25;
reg[15:0] r_22_26;
reg[15:0] r_22_27;
reg[15:0] r_22_28;
reg[15:0] r_22_29;
reg[15:0] r_22_30;
reg[15:0] r_22_31;
reg[15:0] r_22_32;
reg[15:0] r_22_33;
reg[15:0] r_22_34;
reg[15:0] r_22_35;
reg[15:0] r_22_36;
reg[15:0] r_22_37;
reg[15:0] r_22_38;
reg[15:0] r_22_39;
reg[15:0] r_22_40;
reg[15:0] r_22_41;
reg[15:0] r_22_42;
reg[15:0] r_22_43;
reg[15:0] r_22_44;
reg[15:0] r_22_45;
reg[15:0] r_22_46;
reg[15:0] r_22_47;
reg[15:0] r_22_48;
reg[15:0] r_22_49;
reg[15:0] r_22_50;
reg[15:0] r_22_51;
reg[15:0] r_22_52;
reg[15:0] r_22_53;
reg[15:0] r_22_54;
reg[15:0] r_22_55;
reg[15:0] r_22_56;
reg[15:0] r_22_57;
reg[15:0] r_22_58;
reg[15:0] r_22_59;
reg[15:0] r_22_60;
reg[15:0] r_22_61;
reg[15:0] r_22_62;
reg[15:0] r_22_63;
reg[15:0] r_23_0;
reg[15:0] r_23_1;
reg[15:0] r_23_2;
reg[15:0] r_23_3;
reg[15:0] r_23_4;
reg[15:0] r_23_5;
reg[15:0] r_23_6;
reg[15:0] r_23_7;
reg[15:0] r_23_8;
reg[15:0] r_23_9;
reg[15:0] r_23_10;
reg[15:0] r_23_11;
reg[15:0] r_23_12;
reg[15:0] r_23_13;
reg[15:0] r_23_14;
reg[15:0] r_23_15;
reg[15:0] r_23_16;
reg[15:0] r_23_17;
reg[15:0] r_23_18;
reg[15:0] r_23_19;
reg[15:0] r_23_20;
reg[15:0] r_23_21;
reg[15:0] r_23_22;
reg[15:0] r_23_23;
reg[15:0] r_23_24;
reg[15:0] r_23_25;
reg[15:0] r_23_26;
reg[15:0] r_23_27;
reg[15:0] r_23_28;
reg[15:0] r_23_29;
reg[15:0] r_23_30;
reg[15:0] r_23_31;
reg[15:0] r_23_32;
reg[15:0] r_23_33;
reg[15:0] r_23_34;
reg[15:0] r_23_35;
reg[15:0] r_23_36;
reg[15:0] r_23_37;
reg[15:0] r_23_38;
reg[15:0] r_23_39;
reg[15:0] r_23_40;
reg[15:0] r_23_41;
reg[15:0] r_23_42;
reg[15:0] r_23_43;
reg[15:0] r_23_44;
reg[15:0] r_23_45;
reg[15:0] r_23_46;
reg[15:0] r_23_47;
reg[15:0] r_23_48;
reg[15:0] r_23_49;
reg[15:0] r_23_50;
reg[15:0] r_23_51;
reg[15:0] r_23_52;
reg[15:0] r_23_53;
reg[15:0] r_23_54;
reg[15:0] r_23_55;
reg[15:0] r_23_56;
reg[15:0] r_23_57;
reg[15:0] r_23_58;
reg[15:0] r_23_59;
reg[15:0] r_23_60;
reg[15:0] r_23_61;
reg[15:0] r_23_62;
reg[15:0] r_23_63;
reg[15:0] r_24_0;
reg[15:0] r_24_1;
reg[15:0] r_24_2;
reg[15:0] r_24_3;
reg[15:0] r_24_4;
reg[15:0] r_24_5;
reg[15:0] r_24_6;
reg[15:0] r_24_7;
reg[15:0] r_24_8;
reg[15:0] r_24_9;
reg[15:0] r_24_10;
reg[15:0] r_24_11;
reg[15:0] r_24_12;
reg[15:0] r_24_13;
reg[15:0] r_24_14;
reg[15:0] r_24_15;
reg[15:0] r_24_16;
reg[15:0] r_24_17;
reg[15:0] r_24_18;
reg[15:0] r_24_19;
reg[15:0] r_24_20;
reg[15:0] r_24_21;
reg[15:0] r_24_22;
reg[15:0] r_24_23;
reg[15:0] r_24_24;
reg[15:0] r_24_25;
reg[15:0] r_24_26;
reg[15:0] r_24_27;
reg[15:0] r_24_28;
reg[15:0] r_24_29;
reg[15:0] r_24_30;
reg[15:0] r_24_31;
reg[15:0] r_24_32;
reg[15:0] r_24_33;
reg[15:0] r_24_34;
reg[15:0] r_24_35;
reg[15:0] r_24_36;
reg[15:0] r_24_37;
reg[15:0] r_24_38;
reg[15:0] r_24_39;
reg[15:0] r_24_40;
reg[15:0] r_24_41;
reg[15:0] r_24_42;
reg[15:0] r_24_43;
reg[15:0] r_24_44;
reg[15:0] r_24_45;
reg[15:0] r_24_46;
reg[15:0] r_24_47;
reg[15:0] r_24_48;
reg[15:0] r_24_49;
reg[15:0] r_24_50;
reg[15:0] r_24_51;
reg[15:0] r_24_52;
reg[15:0] r_24_53;
reg[15:0] r_24_54;
reg[15:0] r_24_55;
reg[15:0] r_24_56;
reg[15:0] r_24_57;
reg[15:0] r_24_58;
reg[15:0] r_24_59;
reg[15:0] r_24_60;
reg[15:0] r_24_61;
reg[15:0] r_24_62;
reg[15:0] r_24_63;
reg[15:0] r_25_0;
reg[15:0] r_25_1;
reg[15:0] r_25_2;
reg[15:0] r_25_3;
reg[15:0] r_25_4;
reg[15:0] r_25_5;
reg[15:0] r_25_6;
reg[15:0] r_25_7;
reg[15:0] r_25_8;
reg[15:0] r_25_9;
reg[15:0] r_25_10;
reg[15:0] r_25_11;
reg[15:0] r_25_12;
reg[15:0] r_25_13;
reg[15:0] r_25_14;
reg[15:0] r_25_15;
reg[15:0] r_25_16;
reg[15:0] r_25_17;
reg[15:0] r_25_18;
reg[15:0] r_25_19;
reg[15:0] r_25_20;
reg[15:0] r_25_21;
reg[15:0] r_25_22;
reg[15:0] r_25_23;
reg[15:0] r_25_24;
reg[15:0] r_25_25;
reg[15:0] r_25_26;
reg[15:0] r_25_27;
reg[15:0] r_25_28;
reg[15:0] r_25_29;
reg[15:0] r_25_30;
reg[15:0] r_25_31;
reg[15:0] r_25_32;
reg[15:0] r_25_33;
reg[15:0] r_25_34;
reg[15:0] r_25_35;
reg[15:0] r_25_36;
reg[15:0] r_25_37;
reg[15:0] r_25_38;
reg[15:0] r_25_39;
reg[15:0] r_25_40;
reg[15:0] r_25_41;
reg[15:0] r_25_42;
reg[15:0] r_25_43;
reg[15:0] r_25_44;
reg[15:0] r_25_45;
reg[15:0] r_25_46;
reg[15:0] r_25_47;
reg[15:0] r_25_48;
reg[15:0] r_25_49;
reg[15:0] r_25_50;
reg[15:0] r_25_51;
reg[15:0] r_25_52;
reg[15:0] r_25_53;
reg[15:0] r_25_54;
reg[15:0] r_25_55;
reg[15:0] r_25_56;
reg[15:0] r_25_57;
reg[15:0] r_25_58;
reg[15:0] r_25_59;
reg[15:0] r_25_60;
reg[15:0] r_25_61;
reg[15:0] r_25_62;
reg[15:0] r_25_63;
reg[15:0] r_26_0;
reg[15:0] r_26_1;
reg[15:0] r_26_2;
reg[15:0] r_26_3;
reg[15:0] r_26_4;
reg[15:0] r_26_5;
reg[15:0] r_26_6;
reg[15:0] r_26_7;
reg[15:0] r_26_8;
reg[15:0] r_26_9;
reg[15:0] r_26_10;
reg[15:0] r_26_11;
reg[15:0] r_26_12;
reg[15:0] r_26_13;
reg[15:0] r_26_14;
reg[15:0] r_26_15;
reg[15:0] r_26_16;
reg[15:0] r_26_17;
reg[15:0] r_26_18;
reg[15:0] r_26_19;
reg[15:0] r_26_20;
reg[15:0] r_26_21;
reg[15:0] r_26_22;
reg[15:0] r_26_23;
reg[15:0] r_26_24;
reg[15:0] r_26_25;
reg[15:0] r_26_26;
reg[15:0] r_26_27;
reg[15:0] r_26_28;
reg[15:0] r_26_29;
reg[15:0] r_26_30;
reg[15:0] r_26_31;
reg[15:0] r_26_32;
reg[15:0] r_26_33;
reg[15:0] r_26_34;
reg[15:0] r_26_35;
reg[15:0] r_26_36;
reg[15:0] r_26_37;
reg[15:0] r_26_38;
reg[15:0] r_26_39;
reg[15:0] r_26_40;
reg[15:0] r_26_41;
reg[15:0] r_26_42;
reg[15:0] r_26_43;
reg[15:0] r_26_44;
reg[15:0] r_26_45;
reg[15:0] r_26_46;
reg[15:0] r_26_47;
reg[15:0] r_26_48;
reg[15:0] r_26_49;
reg[15:0] r_26_50;
reg[15:0] r_26_51;
reg[15:0] r_26_52;
reg[15:0] r_26_53;
reg[15:0] r_26_54;
reg[15:0] r_26_55;
reg[15:0] r_26_56;
reg[15:0] r_26_57;
reg[15:0] r_26_58;
reg[15:0] r_26_59;
reg[15:0] r_26_60;
reg[15:0] r_26_61;
reg[15:0] r_26_62;
reg[15:0] r_26_63;
reg[15:0] r_27_0;
reg[15:0] r_27_1;
reg[15:0] r_27_2;
reg[15:0] r_27_3;
reg[15:0] r_27_4;
reg[15:0] r_27_5;
reg[15:0] r_27_6;
reg[15:0] r_27_7;
reg[15:0] r_27_8;
reg[15:0] r_27_9;
reg[15:0] r_27_10;
reg[15:0] r_27_11;
reg[15:0] r_27_12;
reg[15:0] r_27_13;
reg[15:0] r_27_14;
reg[15:0] r_27_15;
reg[15:0] r_27_16;
reg[15:0] r_27_17;
reg[15:0] r_27_18;
reg[15:0] r_27_19;
reg[15:0] r_27_20;
reg[15:0] r_27_21;
reg[15:0] r_27_22;
reg[15:0] r_27_23;
reg[15:0] r_27_24;
reg[15:0] r_27_25;
reg[15:0] r_27_26;
reg[15:0] r_27_27;
reg[15:0] r_27_28;
reg[15:0] r_27_29;
reg[15:0] r_27_30;
reg[15:0] r_27_31;
reg[15:0] r_27_32;
reg[15:0] r_27_33;
reg[15:0] r_27_34;
reg[15:0] r_27_35;
reg[15:0] r_27_36;
reg[15:0] r_27_37;
reg[15:0] r_27_38;
reg[15:0] r_27_39;
reg[15:0] r_27_40;
reg[15:0] r_27_41;
reg[15:0] r_27_42;
reg[15:0] r_27_43;
reg[15:0] r_27_44;
reg[15:0] r_27_45;
reg[15:0] r_27_46;
reg[15:0] r_27_47;
reg[15:0] r_27_48;
reg[15:0] r_27_49;
reg[15:0] r_27_50;
reg[15:0] r_27_51;
reg[15:0] r_27_52;
reg[15:0] r_27_53;
reg[15:0] r_27_54;
reg[15:0] r_27_55;
reg[15:0] r_27_56;
reg[15:0] r_27_57;
reg[15:0] r_27_58;
reg[15:0] r_27_59;
reg[15:0] r_27_60;
reg[15:0] r_27_61;
reg[15:0] r_27_62;
reg[15:0] r_27_63;
reg[15:0] r_28_0;
reg[15:0] r_28_1;
reg[15:0] r_28_2;
reg[15:0] r_28_3;
reg[15:0] r_28_4;
reg[15:0] r_28_5;
reg[15:0] r_28_6;
reg[15:0] r_28_7;
reg[15:0] r_28_8;
reg[15:0] r_28_9;
reg[15:0] r_28_10;
reg[15:0] r_28_11;
reg[15:0] r_28_12;
reg[15:0] r_28_13;
reg[15:0] r_28_14;
reg[15:0] r_28_15;
reg[15:0] r_28_16;
reg[15:0] r_28_17;
reg[15:0] r_28_18;
reg[15:0] r_28_19;
reg[15:0] r_28_20;
reg[15:0] r_28_21;
reg[15:0] r_28_22;
reg[15:0] r_28_23;
reg[15:0] r_28_24;
reg[15:0] r_28_25;
reg[15:0] r_28_26;
reg[15:0] r_28_27;
reg[15:0] r_28_28;
reg[15:0] r_28_29;
reg[15:0] r_28_30;
reg[15:0] r_28_31;
reg[15:0] r_28_32;
reg[15:0] r_28_33;
reg[15:0] r_28_34;
reg[15:0] r_28_35;
reg[15:0] r_28_36;
reg[15:0] r_28_37;
reg[15:0] r_28_38;
reg[15:0] r_28_39;
reg[15:0] r_28_40;
reg[15:0] r_28_41;
reg[15:0] r_28_42;
reg[15:0] r_28_43;
reg[15:0] r_28_44;
reg[15:0] r_28_45;
reg[15:0] r_28_46;
reg[15:0] r_28_47;
reg[15:0] r_28_48;
reg[15:0] r_28_49;
reg[15:0] r_28_50;
reg[15:0] r_28_51;
reg[15:0] r_28_52;
reg[15:0] r_28_53;
reg[15:0] r_28_54;
reg[15:0] r_28_55;
reg[15:0] r_28_56;
reg[15:0] r_28_57;
reg[15:0] r_28_58;
reg[15:0] r_28_59;
reg[15:0] r_28_60;
reg[15:0] r_28_61;
reg[15:0] r_28_62;
reg[15:0] r_28_63;
reg[15:0] r_29_0;
reg[15:0] r_29_1;
reg[15:0] r_29_2;
reg[15:0] r_29_3;
reg[15:0] r_29_4;
reg[15:0] r_29_5;
reg[15:0] r_29_6;
reg[15:0] r_29_7;
reg[15:0] r_29_8;
reg[15:0] r_29_9;
reg[15:0] r_29_10;
reg[15:0] r_29_11;
reg[15:0] r_29_12;
reg[15:0] r_29_13;
reg[15:0] r_29_14;
reg[15:0] r_29_15;
reg[15:0] r_29_16;
reg[15:0] r_29_17;
reg[15:0] r_29_18;
reg[15:0] r_29_19;
reg[15:0] r_29_20;
reg[15:0] r_29_21;
reg[15:0] r_29_22;
reg[15:0] r_29_23;
reg[15:0] r_29_24;
reg[15:0] r_29_25;
reg[15:0] r_29_26;
reg[15:0] r_29_27;
reg[15:0] r_29_28;
reg[15:0] r_29_29;
reg[15:0] r_29_30;
reg[15:0] r_29_31;
reg[15:0] r_29_32;
reg[15:0] r_29_33;
reg[15:0] r_29_34;
reg[15:0] r_29_35;
reg[15:0] r_29_36;
reg[15:0] r_29_37;
reg[15:0] r_29_38;
reg[15:0] r_29_39;
reg[15:0] r_29_40;
reg[15:0] r_29_41;
reg[15:0] r_29_42;
reg[15:0] r_29_43;
reg[15:0] r_29_44;
reg[15:0] r_29_45;
reg[15:0] r_29_46;
reg[15:0] r_29_47;
reg[15:0] r_29_48;
reg[15:0] r_29_49;
reg[15:0] r_29_50;
reg[15:0] r_29_51;
reg[15:0] r_29_52;
reg[15:0] r_29_53;
reg[15:0] r_29_54;
reg[15:0] r_29_55;
reg[15:0] r_29_56;
reg[15:0] r_29_57;
reg[15:0] r_29_58;
reg[15:0] r_29_59;
reg[15:0] r_29_60;
reg[15:0] r_29_61;
reg[15:0] r_29_62;
reg[15:0] r_29_63;
reg[15:0] r_30_0;
reg[15:0] r_30_1;
reg[15:0] r_30_2;
reg[15:0] r_30_3;
reg[15:0] r_30_4;
reg[15:0] r_30_5;
reg[15:0] r_30_6;
reg[15:0] r_30_7;
reg[15:0] r_30_8;
reg[15:0] r_30_9;
reg[15:0] r_30_10;
reg[15:0] r_30_11;
reg[15:0] r_30_12;
reg[15:0] r_30_13;
reg[15:0] r_30_14;
reg[15:0] r_30_15;
reg[15:0] r_30_16;
reg[15:0] r_30_17;
reg[15:0] r_30_18;
reg[15:0] r_30_19;
reg[15:0] r_30_20;
reg[15:0] r_30_21;
reg[15:0] r_30_22;
reg[15:0] r_30_23;
reg[15:0] r_30_24;
reg[15:0] r_30_25;
reg[15:0] r_30_26;
reg[15:0] r_30_27;
reg[15:0] r_30_28;
reg[15:0] r_30_29;
reg[15:0] r_30_30;
reg[15:0] r_30_31;
reg[15:0] r_30_32;
reg[15:0] r_30_33;
reg[15:0] r_30_34;
reg[15:0] r_30_35;
reg[15:0] r_30_36;
reg[15:0] r_30_37;
reg[15:0] r_30_38;
reg[15:0] r_30_39;
reg[15:0] r_30_40;
reg[15:0] r_30_41;
reg[15:0] r_30_42;
reg[15:0] r_30_43;
reg[15:0] r_30_44;
reg[15:0] r_30_45;
reg[15:0] r_30_46;
reg[15:0] r_30_47;
reg[15:0] r_30_48;
reg[15:0] r_30_49;
reg[15:0] r_30_50;
reg[15:0] r_30_51;
reg[15:0] r_30_52;
reg[15:0] r_30_53;
reg[15:0] r_30_54;
reg[15:0] r_30_55;
reg[15:0] r_30_56;
reg[15:0] r_30_57;
reg[15:0] r_30_58;
reg[15:0] r_30_59;
reg[15:0] r_30_60;
reg[15:0] r_30_61;
reg[15:0] r_30_62;
reg[15:0] r_30_63;
reg[15:0] r_31_0;
reg[15:0] r_31_1;
reg[15:0] r_31_2;
reg[15:0] r_31_3;
reg[15:0] r_31_4;
reg[15:0] r_31_5;
reg[15:0] r_31_6;
reg[15:0] r_31_7;
reg[15:0] r_31_8;
reg[15:0] r_31_9;
reg[15:0] r_31_10;
reg[15:0] r_31_11;
reg[15:0] r_31_12;
reg[15:0] r_31_13;
reg[15:0] r_31_14;
reg[15:0] r_31_15;
reg[15:0] r_31_16;
reg[15:0] r_31_17;
reg[15:0] r_31_18;
reg[15:0] r_31_19;
reg[15:0] r_31_20;
reg[15:0] r_31_21;
reg[15:0] r_31_22;
reg[15:0] r_31_23;
reg[15:0] r_31_24;
reg[15:0] r_31_25;
reg[15:0] r_31_26;
reg[15:0] r_31_27;
reg[15:0] r_31_28;
reg[15:0] r_31_29;
reg[15:0] r_31_30;
reg[15:0] r_31_31;
reg[15:0] r_31_32;
reg[15:0] r_31_33;
reg[15:0] r_31_34;
reg[15:0] r_31_35;
reg[15:0] r_31_36;
reg[15:0] r_31_37;
reg[15:0] r_31_38;
reg[15:0] r_31_39;
reg[15:0] r_31_40;
reg[15:0] r_31_41;
reg[15:0] r_31_42;
reg[15:0] r_31_43;
reg[15:0] r_31_44;
reg[15:0] r_31_45;
reg[15:0] r_31_46;
reg[15:0] r_31_47;
reg[15:0] r_31_48;
reg[15:0] r_31_49;
reg[15:0] r_31_50;
reg[15:0] r_31_51;
reg[15:0] r_31_52;
reg[15:0] r_31_53;
reg[15:0] r_31_54;
reg[15:0] r_31_55;
reg[15:0] r_31_56;
reg[15:0] r_31_57;
reg[15:0] r_31_58;
reg[15:0] r_31_59;
reg[15:0] r_31_60;
reg[15:0] r_31_61;
reg[15:0] r_31_62;
reg[15:0] r_31_63;
reg[15:0] r_32_0;
reg[15:0] r_32_1;
reg[15:0] r_32_2;
reg[15:0] r_32_3;
reg[15:0] r_32_4;
reg[15:0] r_32_5;
reg[15:0] r_32_6;
reg[15:0] r_32_7;
reg[15:0] r_32_8;
reg[15:0] r_32_9;
reg[15:0] r_32_10;
reg[15:0] r_32_11;
reg[15:0] r_32_12;
reg[15:0] r_32_13;
reg[15:0] r_32_14;
reg[15:0] r_32_15;
reg[15:0] r_32_16;
reg[15:0] r_32_17;
reg[15:0] r_32_18;
reg[15:0] r_32_19;
reg[15:0] r_32_20;
reg[15:0] r_32_21;
reg[15:0] r_32_22;
reg[15:0] r_32_23;
reg[15:0] r_32_24;
reg[15:0] r_32_25;
reg[15:0] r_32_26;
reg[15:0] r_32_27;
reg[15:0] r_32_28;
reg[15:0] r_32_29;
reg[15:0] r_32_30;
reg[15:0] r_32_31;
reg[15:0] r_32_32;
reg[15:0] r_32_33;
reg[15:0] r_32_34;
reg[15:0] r_32_35;
reg[15:0] r_32_36;
reg[15:0] r_32_37;
reg[15:0] r_32_38;
reg[15:0] r_32_39;
reg[15:0] r_32_40;
reg[15:0] r_32_41;
reg[15:0] r_32_42;
reg[15:0] r_32_43;
reg[15:0] r_32_44;
reg[15:0] r_32_45;
reg[15:0] r_32_46;
reg[15:0] r_32_47;
reg[15:0] r_32_48;
reg[15:0] r_32_49;
reg[15:0] r_32_50;
reg[15:0] r_32_51;
reg[15:0] r_32_52;
reg[15:0] r_32_53;
reg[15:0] r_32_54;
reg[15:0] r_32_55;
reg[15:0] r_32_56;
reg[15:0] r_32_57;
reg[15:0] r_32_58;
reg[15:0] r_32_59;
reg[15:0] r_32_60;
reg[15:0] r_32_61;
reg[15:0] r_32_62;
reg[15:0] r_32_63;
reg[15:0] r_33_0;
reg[15:0] r_33_1;
reg[15:0] r_33_2;
reg[15:0] r_33_3;
reg[15:0] r_33_4;
reg[15:0] r_33_5;
reg[15:0] r_33_6;
reg[15:0] r_33_7;
reg[15:0] r_33_8;
reg[15:0] r_33_9;
reg[15:0] r_33_10;
reg[15:0] r_33_11;
reg[15:0] r_33_12;
reg[15:0] r_33_13;
reg[15:0] r_33_14;
reg[15:0] r_33_15;
reg[15:0] r_33_16;
reg[15:0] r_33_17;
reg[15:0] r_33_18;
reg[15:0] r_33_19;
reg[15:0] r_33_20;
reg[15:0] r_33_21;
reg[15:0] r_33_22;
reg[15:0] r_33_23;
reg[15:0] r_33_24;
reg[15:0] r_33_25;
reg[15:0] r_33_26;
reg[15:0] r_33_27;
reg[15:0] r_33_28;
reg[15:0] r_33_29;
reg[15:0] r_33_30;
reg[15:0] r_33_31;
reg[15:0] r_33_32;
reg[15:0] r_33_33;
reg[15:0] r_33_34;
reg[15:0] r_33_35;
reg[15:0] r_33_36;
reg[15:0] r_33_37;
reg[15:0] r_33_38;
reg[15:0] r_33_39;
reg[15:0] r_33_40;
reg[15:0] r_33_41;
reg[15:0] r_33_42;
reg[15:0] r_33_43;
reg[15:0] r_33_44;
reg[15:0] r_33_45;
reg[15:0] r_33_46;
reg[15:0] r_33_47;
reg[15:0] r_33_48;
reg[15:0] r_33_49;
reg[15:0] r_33_50;
reg[15:0] r_33_51;
reg[15:0] r_33_52;
reg[15:0] r_33_53;
reg[15:0] r_33_54;
reg[15:0] r_33_55;
reg[15:0] r_33_56;
reg[15:0] r_33_57;
reg[15:0] r_33_58;
reg[15:0] r_33_59;
reg[15:0] r_33_60;
reg[15:0] r_33_61;
reg[15:0] r_33_62;
reg[15:0] r_33_63;
reg[15:0] r_34_0;
reg[15:0] r_34_1;
reg[15:0] r_34_2;
reg[15:0] r_34_3;
reg[15:0] r_34_4;
reg[15:0] r_34_5;
reg[15:0] r_34_6;
reg[15:0] r_34_7;
reg[15:0] r_34_8;
reg[15:0] r_34_9;
reg[15:0] r_34_10;
reg[15:0] r_34_11;
reg[15:0] r_34_12;
reg[15:0] r_34_13;
reg[15:0] r_34_14;
reg[15:0] r_34_15;
reg[15:0] r_34_16;
reg[15:0] r_34_17;
reg[15:0] r_34_18;
reg[15:0] r_34_19;
reg[15:0] r_34_20;
reg[15:0] r_34_21;
reg[15:0] r_34_22;
reg[15:0] r_34_23;
reg[15:0] r_34_24;
reg[15:0] r_34_25;
reg[15:0] r_34_26;
reg[15:0] r_34_27;
reg[15:0] r_34_28;
reg[15:0] r_34_29;
reg[15:0] r_34_30;
reg[15:0] r_34_31;
reg[15:0] r_34_32;
reg[15:0] r_34_33;
reg[15:0] r_34_34;
reg[15:0] r_34_35;
reg[15:0] r_34_36;
reg[15:0] r_34_37;
reg[15:0] r_34_38;
reg[15:0] r_34_39;
reg[15:0] r_34_40;
reg[15:0] r_34_41;
reg[15:0] r_34_42;
reg[15:0] r_34_43;
reg[15:0] r_34_44;
reg[15:0] r_34_45;
reg[15:0] r_34_46;
reg[15:0] r_34_47;
reg[15:0] r_34_48;
reg[15:0] r_34_49;
reg[15:0] r_34_50;
reg[15:0] r_34_51;
reg[15:0] r_34_52;
reg[15:0] r_34_53;
reg[15:0] r_34_54;
reg[15:0] r_34_55;
reg[15:0] r_34_56;
reg[15:0] r_34_57;
reg[15:0] r_34_58;
reg[15:0] r_34_59;
reg[15:0] r_34_60;
reg[15:0] r_34_61;
reg[15:0] r_34_62;
reg[15:0] r_34_63;
reg[15:0] r_35_0;
reg[15:0] r_35_1;
reg[15:0] r_35_2;
reg[15:0] r_35_3;
reg[15:0] r_35_4;
reg[15:0] r_35_5;
reg[15:0] r_35_6;
reg[15:0] r_35_7;
reg[15:0] r_35_8;
reg[15:0] r_35_9;
reg[15:0] r_35_10;
reg[15:0] r_35_11;
reg[15:0] r_35_12;
reg[15:0] r_35_13;
reg[15:0] r_35_14;
reg[15:0] r_35_15;
reg[15:0] r_35_16;
reg[15:0] r_35_17;
reg[15:0] r_35_18;
reg[15:0] r_35_19;
reg[15:0] r_35_20;
reg[15:0] r_35_21;
reg[15:0] r_35_22;
reg[15:0] r_35_23;
reg[15:0] r_35_24;
reg[15:0] r_35_25;
reg[15:0] r_35_26;
reg[15:0] r_35_27;
reg[15:0] r_35_28;
reg[15:0] r_35_29;
reg[15:0] r_35_30;
reg[15:0] r_35_31;
reg[15:0] r_35_32;
reg[15:0] r_35_33;
reg[15:0] r_35_34;
reg[15:0] r_35_35;
reg[15:0] r_35_36;
reg[15:0] r_35_37;
reg[15:0] r_35_38;
reg[15:0] r_35_39;
reg[15:0] r_35_40;
reg[15:0] r_35_41;
reg[15:0] r_35_42;
reg[15:0] r_35_43;
reg[15:0] r_35_44;
reg[15:0] r_35_45;
reg[15:0] r_35_46;
reg[15:0] r_35_47;
reg[15:0] r_35_48;
reg[15:0] r_35_49;
reg[15:0] r_35_50;
reg[15:0] r_35_51;
reg[15:0] r_35_52;
reg[15:0] r_35_53;
reg[15:0] r_35_54;
reg[15:0] r_35_55;
reg[15:0] r_35_56;
reg[15:0] r_35_57;
reg[15:0] r_35_58;
reg[15:0] r_35_59;
reg[15:0] r_35_60;
reg[15:0] r_35_61;
reg[15:0] r_35_62;
reg[15:0] r_35_63;
reg[15:0] r_36_0;
reg[15:0] r_36_1;
reg[15:0] r_36_2;
reg[15:0] r_36_3;
reg[15:0] r_36_4;
reg[15:0] r_36_5;
reg[15:0] r_36_6;
reg[15:0] r_36_7;
reg[15:0] r_36_8;
reg[15:0] r_36_9;
reg[15:0] r_36_10;
reg[15:0] r_36_11;
reg[15:0] r_36_12;
reg[15:0] r_36_13;
reg[15:0] r_36_14;
reg[15:0] r_36_15;
reg[15:0] r_36_16;
reg[15:0] r_36_17;
reg[15:0] r_36_18;
reg[15:0] r_36_19;
reg[15:0] r_36_20;
reg[15:0] r_36_21;
reg[15:0] r_36_22;
reg[15:0] r_36_23;
reg[15:0] r_36_24;
reg[15:0] r_36_25;
reg[15:0] r_36_26;
reg[15:0] r_36_27;
reg[15:0] r_36_28;
reg[15:0] r_36_29;
reg[15:0] r_36_30;
reg[15:0] r_36_31;
reg[15:0] r_36_32;
reg[15:0] r_36_33;
reg[15:0] r_36_34;
reg[15:0] r_36_35;
reg[15:0] r_36_36;
reg[15:0] r_36_37;
reg[15:0] r_36_38;
reg[15:0] r_36_39;
reg[15:0] r_36_40;
reg[15:0] r_36_41;
reg[15:0] r_36_42;
reg[15:0] r_36_43;
reg[15:0] r_36_44;
reg[15:0] r_36_45;
reg[15:0] r_36_46;
reg[15:0] r_36_47;
reg[15:0] r_36_48;
reg[15:0] r_36_49;
reg[15:0] r_36_50;
reg[15:0] r_36_51;
reg[15:0] r_36_52;
reg[15:0] r_36_53;
reg[15:0] r_36_54;
reg[15:0] r_36_55;
reg[15:0] r_36_56;
reg[15:0] r_36_57;
reg[15:0] r_36_58;
reg[15:0] r_36_59;
reg[15:0] r_36_60;
reg[15:0] r_36_61;
reg[15:0] r_36_62;
reg[15:0] r_36_63;
reg[15:0] r_37_0;
reg[15:0] r_37_1;
reg[15:0] r_37_2;
reg[15:0] r_37_3;
reg[15:0] r_37_4;
reg[15:0] r_37_5;
reg[15:0] r_37_6;
reg[15:0] r_37_7;
reg[15:0] r_37_8;
reg[15:0] r_37_9;
reg[15:0] r_37_10;
reg[15:0] r_37_11;
reg[15:0] r_37_12;
reg[15:0] r_37_13;
reg[15:0] r_37_14;
reg[15:0] r_37_15;
reg[15:0] r_37_16;
reg[15:0] r_37_17;
reg[15:0] r_37_18;
reg[15:0] r_37_19;
reg[15:0] r_37_20;
reg[15:0] r_37_21;
reg[15:0] r_37_22;
reg[15:0] r_37_23;
reg[15:0] r_37_24;
reg[15:0] r_37_25;
reg[15:0] r_37_26;
reg[15:0] r_37_27;
reg[15:0] r_37_28;
reg[15:0] r_37_29;
reg[15:0] r_37_30;
reg[15:0] r_37_31;
reg[15:0] r_37_32;
reg[15:0] r_37_33;
reg[15:0] r_37_34;
reg[15:0] r_37_35;
reg[15:0] r_37_36;
reg[15:0] r_37_37;
reg[15:0] r_37_38;
reg[15:0] r_37_39;
reg[15:0] r_37_40;
reg[15:0] r_37_41;
reg[15:0] r_37_42;
reg[15:0] r_37_43;
reg[15:0] r_37_44;
reg[15:0] r_37_45;
reg[15:0] r_37_46;
reg[15:0] r_37_47;
reg[15:0] r_37_48;
reg[15:0] r_37_49;
reg[15:0] r_37_50;
reg[15:0] r_37_51;
reg[15:0] r_37_52;
reg[15:0] r_37_53;
reg[15:0] r_37_54;
reg[15:0] r_37_55;
reg[15:0] r_37_56;
reg[15:0] r_37_57;
reg[15:0] r_37_58;
reg[15:0] r_37_59;
reg[15:0] r_37_60;
reg[15:0] r_37_61;
reg[15:0] r_37_62;
reg[15:0] r_37_63;
reg[15:0] r_38_0;
reg[15:0] r_38_1;
reg[15:0] r_38_2;
reg[15:0] r_38_3;
reg[15:0] r_38_4;
reg[15:0] r_38_5;
reg[15:0] r_38_6;
reg[15:0] r_38_7;
reg[15:0] r_38_8;
reg[15:0] r_38_9;
reg[15:0] r_38_10;
reg[15:0] r_38_11;
reg[15:0] r_38_12;
reg[15:0] r_38_13;
reg[15:0] r_38_14;
reg[15:0] r_38_15;
reg[15:0] r_38_16;
reg[15:0] r_38_17;
reg[15:0] r_38_18;
reg[15:0] r_38_19;
reg[15:0] r_38_20;
reg[15:0] r_38_21;
reg[15:0] r_38_22;
reg[15:0] r_38_23;
reg[15:0] r_38_24;
reg[15:0] r_38_25;
reg[15:0] r_38_26;
reg[15:0] r_38_27;
reg[15:0] r_38_28;
reg[15:0] r_38_29;
reg[15:0] r_38_30;
reg[15:0] r_38_31;
reg[15:0] r_38_32;
reg[15:0] r_38_33;
reg[15:0] r_38_34;
reg[15:0] r_38_35;
reg[15:0] r_38_36;
reg[15:0] r_38_37;
reg[15:0] r_38_38;
reg[15:0] r_38_39;
reg[15:0] r_38_40;
reg[15:0] r_38_41;
reg[15:0] r_38_42;
reg[15:0] r_38_43;
reg[15:0] r_38_44;
reg[15:0] r_38_45;
reg[15:0] r_38_46;
reg[15:0] r_38_47;
reg[15:0] r_38_48;
reg[15:0] r_38_49;
reg[15:0] r_38_50;
reg[15:0] r_38_51;
reg[15:0] r_38_52;
reg[15:0] r_38_53;
reg[15:0] r_38_54;
reg[15:0] r_38_55;
reg[15:0] r_38_56;
reg[15:0] r_38_57;
reg[15:0] r_38_58;
reg[15:0] r_38_59;
reg[15:0] r_38_60;
reg[15:0] r_38_61;
reg[15:0] r_38_62;
reg[15:0] r_38_63;
reg[15:0] r_39_0;
reg[15:0] r_39_1;
reg[15:0] r_39_2;
reg[15:0] r_39_3;
reg[15:0] r_39_4;
reg[15:0] r_39_5;
reg[15:0] r_39_6;
reg[15:0] r_39_7;
reg[15:0] r_39_8;
reg[15:0] r_39_9;
reg[15:0] r_39_10;
reg[15:0] r_39_11;
reg[15:0] r_39_12;
reg[15:0] r_39_13;
reg[15:0] r_39_14;
reg[15:0] r_39_15;
reg[15:0] r_39_16;
reg[15:0] r_39_17;
reg[15:0] r_39_18;
reg[15:0] r_39_19;
reg[15:0] r_39_20;
reg[15:0] r_39_21;
reg[15:0] r_39_22;
reg[15:0] r_39_23;
reg[15:0] r_39_24;
reg[15:0] r_39_25;
reg[15:0] r_39_26;
reg[15:0] r_39_27;
reg[15:0] r_39_28;
reg[15:0] r_39_29;
reg[15:0] r_39_30;
reg[15:0] r_39_31;
reg[15:0] r_39_32;
reg[15:0] r_39_33;
reg[15:0] r_39_34;
reg[15:0] r_39_35;
reg[15:0] r_39_36;
reg[15:0] r_39_37;
reg[15:0] r_39_38;
reg[15:0] r_39_39;
reg[15:0] r_39_40;
reg[15:0] r_39_41;
reg[15:0] r_39_42;
reg[15:0] r_39_43;
reg[15:0] r_39_44;
reg[15:0] r_39_45;
reg[15:0] r_39_46;
reg[15:0] r_39_47;
reg[15:0] r_39_48;
reg[15:0] r_39_49;
reg[15:0] r_39_50;
reg[15:0] r_39_51;
reg[15:0] r_39_52;
reg[15:0] r_39_53;
reg[15:0] r_39_54;
reg[15:0] r_39_55;
reg[15:0] r_39_56;
reg[15:0] r_39_57;
reg[15:0] r_39_58;
reg[15:0] r_39_59;
reg[15:0] r_39_60;
reg[15:0] r_39_61;
reg[15:0] r_39_62;
reg[15:0] r_39_63;
reg[15:0] r_40_0;
reg[15:0] r_40_1;
reg[15:0] r_40_2;
reg[15:0] r_40_3;
reg[15:0] r_40_4;
reg[15:0] r_40_5;
reg[15:0] r_40_6;
reg[15:0] r_40_7;
reg[15:0] r_40_8;
reg[15:0] r_40_9;
reg[15:0] r_40_10;
reg[15:0] r_40_11;
reg[15:0] r_40_12;
reg[15:0] r_40_13;
reg[15:0] r_40_14;
reg[15:0] r_40_15;
reg[15:0] r_40_16;
reg[15:0] r_40_17;
reg[15:0] r_40_18;
reg[15:0] r_40_19;
reg[15:0] r_40_20;
reg[15:0] r_40_21;
reg[15:0] r_40_22;
reg[15:0] r_40_23;
reg[15:0] r_40_24;
reg[15:0] r_40_25;
reg[15:0] r_40_26;
reg[15:0] r_40_27;
reg[15:0] r_40_28;
reg[15:0] r_40_29;
reg[15:0] r_40_30;
reg[15:0] r_40_31;
reg[15:0] r_40_32;
reg[15:0] r_40_33;
reg[15:0] r_40_34;
reg[15:0] r_40_35;
reg[15:0] r_40_36;
reg[15:0] r_40_37;
reg[15:0] r_40_38;
reg[15:0] r_40_39;
reg[15:0] r_40_40;
reg[15:0] r_40_41;
reg[15:0] r_40_42;
reg[15:0] r_40_43;
reg[15:0] r_40_44;
reg[15:0] r_40_45;
reg[15:0] r_40_46;
reg[15:0] r_40_47;
reg[15:0] r_40_48;
reg[15:0] r_40_49;
reg[15:0] r_40_50;
reg[15:0] r_40_51;
reg[15:0] r_40_52;
reg[15:0] r_40_53;
reg[15:0] r_40_54;
reg[15:0] r_40_55;
reg[15:0] r_40_56;
reg[15:0] r_40_57;
reg[15:0] r_40_58;
reg[15:0] r_40_59;
reg[15:0] r_40_60;
reg[15:0] r_40_61;
reg[15:0] r_40_62;
reg[15:0] r_40_63;
reg[15:0] r_41_0;
reg[15:0] r_41_1;
reg[15:0] r_41_2;
reg[15:0] r_41_3;
reg[15:0] r_41_4;
reg[15:0] r_41_5;
reg[15:0] r_41_6;
reg[15:0] r_41_7;
reg[15:0] r_41_8;
reg[15:0] r_41_9;
reg[15:0] r_41_10;
reg[15:0] r_41_11;
reg[15:0] r_41_12;
reg[15:0] r_41_13;
reg[15:0] r_41_14;
reg[15:0] r_41_15;
reg[15:0] r_41_16;
reg[15:0] r_41_17;
reg[15:0] r_41_18;
reg[15:0] r_41_19;
reg[15:0] r_41_20;
reg[15:0] r_41_21;
reg[15:0] r_41_22;
reg[15:0] r_41_23;
reg[15:0] r_41_24;
reg[15:0] r_41_25;
reg[15:0] r_41_26;
reg[15:0] r_41_27;
reg[15:0] r_41_28;
reg[15:0] r_41_29;
reg[15:0] r_41_30;
reg[15:0] r_41_31;
reg[15:0] r_41_32;
reg[15:0] r_41_33;
reg[15:0] r_41_34;
reg[15:0] r_41_35;
reg[15:0] r_41_36;
reg[15:0] r_41_37;
reg[15:0] r_41_38;
reg[15:0] r_41_39;
reg[15:0] r_41_40;
reg[15:0] r_41_41;
reg[15:0] r_41_42;
reg[15:0] r_41_43;
reg[15:0] r_41_44;
reg[15:0] r_41_45;
reg[15:0] r_41_46;
reg[15:0] r_41_47;
reg[15:0] r_41_48;
reg[15:0] r_41_49;
reg[15:0] r_41_50;
reg[15:0] r_41_51;
reg[15:0] r_41_52;
reg[15:0] r_41_53;
reg[15:0] r_41_54;
reg[15:0] r_41_55;
reg[15:0] r_41_56;
reg[15:0] r_41_57;
reg[15:0] r_41_58;
reg[15:0] r_41_59;
reg[15:0] r_41_60;
reg[15:0] r_41_61;
reg[15:0] r_41_62;
reg[15:0] r_41_63;
reg[15:0] r_42_0;
reg[15:0] r_42_1;
reg[15:0] r_42_2;
reg[15:0] r_42_3;
reg[15:0] r_42_4;
reg[15:0] r_42_5;
reg[15:0] r_42_6;
reg[15:0] r_42_7;
reg[15:0] r_42_8;
reg[15:0] r_42_9;
reg[15:0] r_42_10;
reg[15:0] r_42_11;
reg[15:0] r_42_12;
reg[15:0] r_42_13;
reg[15:0] r_42_14;
reg[15:0] r_42_15;
reg[15:0] r_42_16;
reg[15:0] r_42_17;
reg[15:0] r_42_18;
reg[15:0] r_42_19;
reg[15:0] r_42_20;
reg[15:0] r_42_21;
reg[15:0] r_42_22;
reg[15:0] r_42_23;
reg[15:0] r_42_24;
reg[15:0] r_42_25;
reg[15:0] r_42_26;
reg[15:0] r_42_27;
reg[15:0] r_42_28;
reg[15:0] r_42_29;
reg[15:0] r_42_30;
reg[15:0] r_42_31;
reg[15:0] r_42_32;
reg[15:0] r_42_33;
reg[15:0] r_42_34;
reg[15:0] r_42_35;
reg[15:0] r_42_36;
reg[15:0] r_42_37;
reg[15:0] r_42_38;
reg[15:0] r_42_39;
reg[15:0] r_42_40;
reg[15:0] r_42_41;
reg[15:0] r_42_42;
reg[15:0] r_42_43;
reg[15:0] r_42_44;
reg[15:0] r_42_45;
reg[15:0] r_42_46;
reg[15:0] r_42_47;
reg[15:0] r_42_48;
reg[15:0] r_42_49;
reg[15:0] r_42_50;
reg[15:0] r_42_51;
reg[15:0] r_42_52;
reg[15:0] r_42_53;
reg[15:0] r_42_54;
reg[15:0] r_42_55;
reg[15:0] r_42_56;
reg[15:0] r_42_57;
reg[15:0] r_42_58;
reg[15:0] r_42_59;
reg[15:0] r_42_60;
reg[15:0] r_42_61;
reg[15:0] r_42_62;
reg[15:0] r_42_63;
reg[15:0] r_43_0;
reg[15:0] r_43_1;
reg[15:0] r_43_2;
reg[15:0] r_43_3;
reg[15:0] r_43_4;
reg[15:0] r_43_5;
reg[15:0] r_43_6;
reg[15:0] r_43_7;
reg[15:0] r_43_8;
reg[15:0] r_43_9;
reg[15:0] r_43_10;
reg[15:0] r_43_11;
reg[15:0] r_43_12;
reg[15:0] r_43_13;
reg[15:0] r_43_14;
reg[15:0] r_43_15;
reg[15:0] r_43_16;
reg[15:0] r_43_17;
reg[15:0] r_43_18;
reg[15:0] r_43_19;
reg[15:0] r_43_20;
reg[15:0] r_43_21;
reg[15:0] r_43_22;
reg[15:0] r_43_23;
reg[15:0] r_43_24;
reg[15:0] r_43_25;
reg[15:0] r_43_26;
reg[15:0] r_43_27;
reg[15:0] r_43_28;
reg[15:0] r_43_29;
reg[15:0] r_43_30;
reg[15:0] r_43_31;
reg[15:0] r_43_32;
reg[15:0] r_43_33;
reg[15:0] r_43_34;
reg[15:0] r_43_35;
reg[15:0] r_43_36;
reg[15:0] r_43_37;
reg[15:0] r_43_38;
reg[15:0] r_43_39;
reg[15:0] r_43_40;
reg[15:0] r_43_41;
reg[15:0] r_43_42;
reg[15:0] r_43_43;
reg[15:0] r_43_44;
reg[15:0] r_43_45;
reg[15:0] r_43_46;
reg[15:0] r_43_47;
reg[15:0] r_43_48;
reg[15:0] r_43_49;
reg[15:0] r_43_50;
reg[15:0] r_43_51;
reg[15:0] r_43_52;
reg[15:0] r_43_53;
reg[15:0] r_43_54;
reg[15:0] r_43_55;
reg[15:0] r_43_56;
reg[15:0] r_43_57;
reg[15:0] r_43_58;
reg[15:0] r_43_59;
reg[15:0] r_43_60;
reg[15:0] r_43_61;
reg[15:0] r_43_62;
reg[15:0] r_43_63;
reg[15:0] r_44_0;
reg[15:0] r_44_1;
reg[15:0] r_44_2;
reg[15:0] r_44_3;
reg[15:0] r_44_4;
reg[15:0] r_44_5;
reg[15:0] r_44_6;
reg[15:0] r_44_7;
reg[15:0] r_44_8;
reg[15:0] r_44_9;
reg[15:0] r_44_10;
reg[15:0] r_44_11;
reg[15:0] r_44_12;
reg[15:0] r_44_13;
reg[15:0] r_44_14;
reg[15:0] r_44_15;
reg[15:0] r_44_16;
reg[15:0] r_44_17;
reg[15:0] r_44_18;
reg[15:0] r_44_19;
reg[15:0] r_44_20;
reg[15:0] r_44_21;
reg[15:0] r_44_22;
reg[15:0] r_44_23;
reg[15:0] r_44_24;
reg[15:0] r_44_25;
reg[15:0] r_44_26;
reg[15:0] r_44_27;
reg[15:0] r_44_28;
reg[15:0] r_44_29;
reg[15:0] r_44_30;
reg[15:0] r_44_31;
reg[15:0] r_44_32;
reg[15:0] r_44_33;
reg[15:0] r_44_34;
reg[15:0] r_44_35;
reg[15:0] r_44_36;
reg[15:0] r_44_37;
reg[15:0] r_44_38;
reg[15:0] r_44_39;
reg[15:0] r_44_40;
reg[15:0] r_44_41;
reg[15:0] r_44_42;
reg[15:0] r_44_43;
reg[15:0] r_44_44;
reg[15:0] r_44_45;
reg[15:0] r_44_46;
reg[15:0] r_44_47;
reg[15:0] r_44_48;
reg[15:0] r_44_49;
reg[15:0] r_44_50;
reg[15:0] r_44_51;
reg[15:0] r_44_52;
reg[15:0] r_44_53;
reg[15:0] r_44_54;
reg[15:0] r_44_55;
reg[15:0] r_44_56;
reg[15:0] r_44_57;
reg[15:0] r_44_58;
reg[15:0] r_44_59;
reg[15:0] r_44_60;
reg[15:0] r_44_61;
reg[15:0] r_44_62;
reg[15:0] r_44_63;
reg[15:0] r_45_0;
reg[15:0] r_45_1;
reg[15:0] r_45_2;
reg[15:0] r_45_3;
reg[15:0] r_45_4;
reg[15:0] r_45_5;
reg[15:0] r_45_6;
reg[15:0] r_45_7;
reg[15:0] r_45_8;
reg[15:0] r_45_9;
reg[15:0] r_45_10;
reg[15:0] r_45_11;
reg[15:0] r_45_12;
reg[15:0] r_45_13;
reg[15:0] r_45_14;
reg[15:0] r_45_15;
reg[15:0] r_45_16;
reg[15:0] r_45_17;
reg[15:0] r_45_18;
reg[15:0] r_45_19;
reg[15:0] r_45_20;
reg[15:0] r_45_21;
reg[15:0] r_45_22;
reg[15:0] r_45_23;
reg[15:0] r_45_24;
reg[15:0] r_45_25;
reg[15:0] r_45_26;
reg[15:0] r_45_27;
reg[15:0] r_45_28;
reg[15:0] r_45_29;
reg[15:0] r_45_30;
reg[15:0] r_45_31;
reg[15:0] r_45_32;
reg[15:0] r_45_33;
reg[15:0] r_45_34;
reg[15:0] r_45_35;
reg[15:0] r_45_36;
reg[15:0] r_45_37;
reg[15:0] r_45_38;
reg[15:0] r_45_39;
reg[15:0] r_45_40;
reg[15:0] r_45_41;
reg[15:0] r_45_42;
reg[15:0] r_45_43;
reg[15:0] r_45_44;
reg[15:0] r_45_45;
reg[15:0] r_45_46;
reg[15:0] r_45_47;
reg[15:0] r_45_48;
reg[15:0] r_45_49;
reg[15:0] r_45_50;
reg[15:0] r_45_51;
reg[15:0] r_45_52;
reg[15:0] r_45_53;
reg[15:0] r_45_54;
reg[15:0] r_45_55;
reg[15:0] r_45_56;
reg[15:0] r_45_57;
reg[15:0] r_45_58;
reg[15:0] r_45_59;
reg[15:0] r_45_60;
reg[15:0] r_45_61;
reg[15:0] r_45_62;
reg[15:0] r_45_63;
reg[15:0] r_46_0;
reg[15:0] r_46_1;
reg[15:0] r_46_2;
reg[15:0] r_46_3;
reg[15:0] r_46_4;
reg[15:0] r_46_5;
reg[15:0] r_46_6;
reg[15:0] r_46_7;
reg[15:0] r_46_8;
reg[15:0] r_46_9;
reg[15:0] r_46_10;
reg[15:0] r_46_11;
reg[15:0] r_46_12;
reg[15:0] r_46_13;
reg[15:0] r_46_14;
reg[15:0] r_46_15;
reg[15:0] r_46_16;
reg[15:0] r_46_17;
reg[15:0] r_46_18;
reg[15:0] r_46_19;
reg[15:0] r_46_20;
reg[15:0] r_46_21;
reg[15:0] r_46_22;
reg[15:0] r_46_23;
reg[15:0] r_46_24;
reg[15:0] r_46_25;
reg[15:0] r_46_26;
reg[15:0] r_46_27;
reg[15:0] r_46_28;
reg[15:0] r_46_29;
reg[15:0] r_46_30;
reg[15:0] r_46_31;
reg[15:0] r_46_32;
reg[15:0] r_46_33;
reg[15:0] r_46_34;
reg[15:0] r_46_35;
reg[15:0] r_46_36;
reg[15:0] r_46_37;
reg[15:0] r_46_38;
reg[15:0] r_46_39;
reg[15:0] r_46_40;
reg[15:0] r_46_41;
reg[15:0] r_46_42;
reg[15:0] r_46_43;
reg[15:0] r_46_44;
reg[15:0] r_46_45;
reg[15:0] r_46_46;
reg[15:0] r_46_47;
reg[15:0] r_46_48;
reg[15:0] r_46_49;
reg[15:0] r_46_50;
reg[15:0] r_46_51;
reg[15:0] r_46_52;
reg[15:0] r_46_53;
reg[15:0] r_46_54;
reg[15:0] r_46_55;
reg[15:0] r_46_56;
reg[15:0] r_46_57;
reg[15:0] r_46_58;
reg[15:0] r_46_59;
reg[15:0] r_46_60;
reg[15:0] r_46_61;
reg[15:0] r_46_62;
reg[15:0] r_46_63;
reg[15:0] r_47_0;
reg[15:0] r_47_1;
reg[15:0] r_47_2;
reg[15:0] r_47_3;
reg[15:0] r_47_4;
reg[15:0] r_47_5;
reg[15:0] r_47_6;
reg[15:0] r_47_7;
reg[15:0] r_47_8;
reg[15:0] r_47_9;
reg[15:0] r_47_10;
reg[15:0] r_47_11;
reg[15:0] r_47_12;
reg[15:0] r_47_13;
reg[15:0] r_47_14;
reg[15:0] r_47_15;
reg[15:0] r_47_16;
reg[15:0] r_47_17;
reg[15:0] r_47_18;
reg[15:0] r_47_19;
reg[15:0] r_47_20;
reg[15:0] r_47_21;
reg[15:0] r_47_22;
reg[15:0] r_47_23;
reg[15:0] r_47_24;
reg[15:0] r_47_25;
reg[15:0] r_47_26;
reg[15:0] r_47_27;
reg[15:0] r_47_28;
reg[15:0] r_47_29;
reg[15:0] r_47_30;
reg[15:0] r_47_31;
reg[15:0] r_47_32;
reg[15:0] r_47_33;
reg[15:0] r_47_34;
reg[15:0] r_47_35;
reg[15:0] r_47_36;
reg[15:0] r_47_37;
reg[15:0] r_47_38;
reg[15:0] r_47_39;
reg[15:0] r_47_40;
reg[15:0] r_47_41;
reg[15:0] r_47_42;
reg[15:0] r_47_43;
reg[15:0] r_47_44;
reg[15:0] r_47_45;
reg[15:0] r_47_46;
reg[15:0] r_47_47;
reg[15:0] r_47_48;
reg[15:0] r_47_49;
reg[15:0] r_47_50;
reg[15:0] r_47_51;
reg[15:0] r_47_52;
reg[15:0] r_47_53;
reg[15:0] r_47_54;
reg[15:0] r_47_55;
reg[15:0] r_47_56;
reg[15:0] r_47_57;
reg[15:0] r_47_58;
reg[15:0] r_47_59;
reg[15:0] r_47_60;
reg[15:0] r_47_61;
reg[15:0] r_47_62;
reg[15:0] r_47_63;
reg[15:0] r_48_0;
reg[15:0] r_48_1;
reg[15:0] r_48_2;
reg[15:0] r_48_3;
reg[15:0] r_48_4;
reg[15:0] r_48_5;
reg[15:0] r_48_6;
reg[15:0] r_48_7;
reg[15:0] r_48_8;
reg[15:0] r_48_9;
reg[15:0] r_48_10;
reg[15:0] r_48_11;
reg[15:0] r_48_12;
reg[15:0] r_48_13;
reg[15:0] r_48_14;
reg[15:0] r_48_15;
reg[15:0] r_48_16;
reg[15:0] r_48_17;
reg[15:0] r_48_18;
reg[15:0] r_48_19;
reg[15:0] r_48_20;
reg[15:0] r_48_21;
reg[15:0] r_48_22;
reg[15:0] r_48_23;
reg[15:0] r_48_24;
reg[15:0] r_48_25;
reg[15:0] r_48_26;
reg[15:0] r_48_27;
reg[15:0] r_48_28;
reg[15:0] r_48_29;
reg[15:0] r_48_30;
reg[15:0] r_48_31;
reg[15:0] r_48_32;
reg[15:0] r_48_33;
reg[15:0] r_48_34;
reg[15:0] r_48_35;
reg[15:0] r_48_36;
reg[15:0] r_48_37;
reg[15:0] r_48_38;
reg[15:0] r_48_39;
reg[15:0] r_48_40;
reg[15:0] r_48_41;
reg[15:0] r_48_42;
reg[15:0] r_48_43;
reg[15:0] r_48_44;
reg[15:0] r_48_45;
reg[15:0] r_48_46;
reg[15:0] r_48_47;
reg[15:0] r_48_48;
reg[15:0] r_48_49;
reg[15:0] r_48_50;
reg[15:0] r_48_51;
reg[15:0] r_48_52;
reg[15:0] r_48_53;
reg[15:0] r_48_54;
reg[15:0] r_48_55;
reg[15:0] r_48_56;
reg[15:0] r_48_57;
reg[15:0] r_48_58;
reg[15:0] r_48_59;
reg[15:0] r_48_60;
reg[15:0] r_48_61;
reg[15:0] r_48_62;
reg[15:0] r_48_63;
reg[15:0] r_49_0;
reg[15:0] r_49_1;
reg[15:0] r_49_2;
reg[15:0] r_49_3;
reg[15:0] r_49_4;
reg[15:0] r_49_5;
reg[15:0] r_49_6;
reg[15:0] r_49_7;
reg[15:0] r_49_8;
reg[15:0] r_49_9;
reg[15:0] r_49_10;
reg[15:0] r_49_11;
reg[15:0] r_49_12;
reg[15:0] r_49_13;
reg[15:0] r_49_14;
reg[15:0] r_49_15;
reg[15:0] r_49_16;
reg[15:0] r_49_17;
reg[15:0] r_49_18;
reg[15:0] r_49_19;
reg[15:0] r_49_20;
reg[15:0] r_49_21;
reg[15:0] r_49_22;
reg[15:0] r_49_23;
reg[15:0] r_49_24;
reg[15:0] r_49_25;
reg[15:0] r_49_26;
reg[15:0] r_49_27;
reg[15:0] r_49_28;
reg[15:0] r_49_29;
reg[15:0] r_49_30;
reg[15:0] r_49_31;
reg[15:0] r_49_32;
reg[15:0] r_49_33;
reg[15:0] r_49_34;
reg[15:0] r_49_35;
reg[15:0] r_49_36;
reg[15:0] r_49_37;
reg[15:0] r_49_38;
reg[15:0] r_49_39;
reg[15:0] r_49_40;
reg[15:0] r_49_41;
reg[15:0] r_49_42;
reg[15:0] r_49_43;
reg[15:0] r_49_44;
reg[15:0] r_49_45;
reg[15:0] r_49_46;
reg[15:0] r_49_47;
reg[15:0] r_49_48;
reg[15:0] r_49_49;
reg[15:0] r_49_50;
reg[15:0] r_49_51;
reg[15:0] r_49_52;
reg[15:0] r_49_53;
reg[15:0] r_49_54;
reg[15:0] r_49_55;
reg[15:0] r_49_56;
reg[15:0] r_49_57;
reg[15:0] r_49_58;
reg[15:0] r_49_59;
reg[15:0] r_49_60;
reg[15:0] r_49_61;
reg[15:0] r_49_62;
reg[15:0] r_49_63;
reg[15:0] r_50_0;
reg[15:0] r_50_1;
reg[15:0] r_50_2;
reg[15:0] r_50_3;
reg[15:0] r_50_4;
reg[15:0] r_50_5;
reg[15:0] r_50_6;
reg[15:0] r_50_7;
reg[15:0] r_50_8;
reg[15:0] r_50_9;
reg[15:0] r_50_10;
reg[15:0] r_50_11;
reg[15:0] r_50_12;
reg[15:0] r_50_13;
reg[15:0] r_50_14;
reg[15:0] r_50_15;
reg[15:0] r_50_16;
reg[15:0] r_50_17;
reg[15:0] r_50_18;
reg[15:0] r_50_19;
reg[15:0] r_50_20;
reg[15:0] r_50_21;
reg[15:0] r_50_22;
reg[15:0] r_50_23;
reg[15:0] r_50_24;
reg[15:0] r_50_25;
reg[15:0] r_50_26;
reg[15:0] r_50_27;
reg[15:0] r_50_28;
reg[15:0] r_50_29;
reg[15:0] r_50_30;
reg[15:0] r_50_31;
reg[15:0] r_50_32;
reg[15:0] r_50_33;
reg[15:0] r_50_34;
reg[15:0] r_50_35;
reg[15:0] r_50_36;
reg[15:0] r_50_37;
reg[15:0] r_50_38;
reg[15:0] r_50_39;
reg[15:0] r_50_40;
reg[15:0] r_50_41;
reg[15:0] r_50_42;
reg[15:0] r_50_43;
reg[15:0] r_50_44;
reg[15:0] r_50_45;
reg[15:0] r_50_46;
reg[15:0] r_50_47;
reg[15:0] r_50_48;
reg[15:0] r_50_49;
reg[15:0] r_50_50;
reg[15:0] r_50_51;
reg[15:0] r_50_52;
reg[15:0] r_50_53;
reg[15:0] r_50_54;
reg[15:0] r_50_55;
reg[15:0] r_50_56;
reg[15:0] r_50_57;
reg[15:0] r_50_58;
reg[15:0] r_50_59;
reg[15:0] r_50_60;
reg[15:0] r_50_61;
reg[15:0] r_50_62;
reg[15:0] r_50_63;
reg[15:0] r_51_0;
reg[15:0] r_51_1;
reg[15:0] r_51_2;
reg[15:0] r_51_3;
reg[15:0] r_51_4;
reg[15:0] r_51_5;
reg[15:0] r_51_6;
reg[15:0] r_51_7;
reg[15:0] r_51_8;
reg[15:0] r_51_9;
reg[15:0] r_51_10;
reg[15:0] r_51_11;
reg[15:0] r_51_12;
reg[15:0] r_51_13;
reg[15:0] r_51_14;
reg[15:0] r_51_15;
reg[15:0] r_51_16;
reg[15:0] r_51_17;
reg[15:0] r_51_18;
reg[15:0] r_51_19;
reg[15:0] r_51_20;
reg[15:0] r_51_21;
reg[15:0] r_51_22;
reg[15:0] r_51_23;
reg[15:0] r_51_24;
reg[15:0] r_51_25;
reg[15:0] r_51_26;
reg[15:0] r_51_27;
reg[15:0] r_51_28;
reg[15:0] r_51_29;
reg[15:0] r_51_30;
reg[15:0] r_51_31;
reg[15:0] r_51_32;
reg[15:0] r_51_33;
reg[15:0] r_51_34;
reg[15:0] r_51_35;
reg[15:0] r_51_36;
reg[15:0] r_51_37;
reg[15:0] r_51_38;
reg[15:0] r_51_39;
reg[15:0] r_51_40;
reg[15:0] r_51_41;
reg[15:0] r_51_42;
reg[15:0] r_51_43;
reg[15:0] r_51_44;
reg[15:0] r_51_45;
reg[15:0] r_51_46;
reg[15:0] r_51_47;
reg[15:0] r_51_48;
reg[15:0] r_51_49;
reg[15:0] r_51_50;
reg[15:0] r_51_51;
reg[15:0] r_51_52;
reg[15:0] r_51_53;
reg[15:0] r_51_54;
reg[15:0] r_51_55;
reg[15:0] r_51_56;
reg[15:0] r_51_57;
reg[15:0] r_51_58;
reg[15:0] r_51_59;
reg[15:0] r_51_60;
reg[15:0] r_51_61;
reg[15:0] r_51_62;
reg[15:0] r_51_63;
reg[15:0] r_52_0;
reg[15:0] r_52_1;
reg[15:0] r_52_2;
reg[15:0] r_52_3;
reg[15:0] r_52_4;
reg[15:0] r_52_5;
reg[15:0] r_52_6;
reg[15:0] r_52_7;
reg[15:0] r_52_8;
reg[15:0] r_52_9;
reg[15:0] r_52_10;
reg[15:0] r_52_11;
reg[15:0] r_52_12;
reg[15:0] r_52_13;
reg[15:0] r_52_14;
reg[15:0] r_52_15;
reg[15:0] r_52_16;
reg[15:0] r_52_17;
reg[15:0] r_52_18;
reg[15:0] r_52_19;
reg[15:0] r_52_20;
reg[15:0] r_52_21;
reg[15:0] r_52_22;
reg[15:0] r_52_23;
reg[15:0] r_52_24;
reg[15:0] r_52_25;
reg[15:0] r_52_26;
reg[15:0] r_52_27;
reg[15:0] r_52_28;
reg[15:0] r_52_29;
reg[15:0] r_52_30;
reg[15:0] r_52_31;
reg[15:0] r_52_32;
reg[15:0] r_52_33;
reg[15:0] r_52_34;
reg[15:0] r_52_35;
reg[15:0] r_52_36;
reg[15:0] r_52_37;
reg[15:0] r_52_38;
reg[15:0] r_52_39;
reg[15:0] r_52_40;
reg[15:0] r_52_41;
reg[15:0] r_52_42;
reg[15:0] r_52_43;
reg[15:0] r_52_44;
reg[15:0] r_52_45;
reg[15:0] r_52_46;
reg[15:0] r_52_47;
reg[15:0] r_52_48;
reg[15:0] r_52_49;
reg[15:0] r_52_50;
reg[15:0] r_52_51;
reg[15:0] r_52_52;
reg[15:0] r_52_53;
reg[15:0] r_52_54;
reg[15:0] r_52_55;
reg[15:0] r_52_56;
reg[15:0] r_52_57;
reg[15:0] r_52_58;
reg[15:0] r_52_59;
reg[15:0] r_52_60;
reg[15:0] r_52_61;
reg[15:0] r_52_62;
reg[15:0] r_52_63;
reg[15:0] r_53_0;
reg[15:0] r_53_1;
reg[15:0] r_53_2;
reg[15:0] r_53_3;
reg[15:0] r_53_4;
reg[15:0] r_53_5;
reg[15:0] r_53_6;
reg[15:0] r_53_7;
reg[15:0] r_53_8;
reg[15:0] r_53_9;
reg[15:0] r_53_10;
reg[15:0] r_53_11;
reg[15:0] r_53_12;
reg[15:0] r_53_13;
reg[15:0] r_53_14;
reg[15:0] r_53_15;
reg[15:0] r_53_16;
reg[15:0] r_53_17;
reg[15:0] r_53_18;
reg[15:0] r_53_19;
reg[15:0] r_53_20;
reg[15:0] r_53_21;
reg[15:0] r_53_22;
reg[15:0] r_53_23;
reg[15:0] r_53_24;
reg[15:0] r_53_25;
reg[15:0] r_53_26;
reg[15:0] r_53_27;
reg[15:0] r_53_28;
reg[15:0] r_53_29;
reg[15:0] r_53_30;
reg[15:0] r_53_31;
reg[15:0] r_53_32;
reg[15:0] r_53_33;
reg[15:0] r_53_34;
reg[15:0] r_53_35;
reg[15:0] r_53_36;
reg[15:0] r_53_37;
reg[15:0] r_53_38;
reg[15:0] r_53_39;
reg[15:0] r_53_40;
reg[15:0] r_53_41;
reg[15:0] r_53_42;
reg[15:0] r_53_43;
reg[15:0] r_53_44;
reg[15:0] r_53_45;
reg[15:0] r_53_46;
reg[15:0] r_53_47;
reg[15:0] r_53_48;
reg[15:0] r_53_49;
reg[15:0] r_53_50;
reg[15:0] r_53_51;
reg[15:0] r_53_52;
reg[15:0] r_53_53;
reg[15:0] r_53_54;
reg[15:0] r_53_55;
reg[15:0] r_53_56;
reg[15:0] r_53_57;
reg[15:0] r_53_58;
reg[15:0] r_53_59;
reg[15:0] r_53_60;
reg[15:0] r_53_61;
reg[15:0] r_53_62;
reg[15:0] r_53_63;
reg[15:0] r_54_0;
reg[15:0] r_54_1;
reg[15:0] r_54_2;
reg[15:0] r_54_3;
reg[15:0] r_54_4;
reg[15:0] r_54_5;
reg[15:0] r_54_6;
reg[15:0] r_54_7;
reg[15:0] r_54_8;
reg[15:0] r_54_9;
reg[15:0] r_54_10;
reg[15:0] r_54_11;
reg[15:0] r_54_12;
reg[15:0] r_54_13;
reg[15:0] r_54_14;
reg[15:0] r_54_15;
reg[15:0] r_54_16;
reg[15:0] r_54_17;
reg[15:0] r_54_18;
reg[15:0] r_54_19;
reg[15:0] r_54_20;
reg[15:0] r_54_21;
reg[15:0] r_54_22;
reg[15:0] r_54_23;
reg[15:0] r_54_24;
reg[15:0] r_54_25;
reg[15:0] r_54_26;
reg[15:0] r_54_27;
reg[15:0] r_54_28;
reg[15:0] r_54_29;
reg[15:0] r_54_30;
reg[15:0] r_54_31;
reg[15:0] r_54_32;
reg[15:0] r_54_33;
reg[15:0] r_54_34;
reg[15:0] r_54_35;
reg[15:0] r_54_36;
reg[15:0] r_54_37;
reg[15:0] r_54_38;
reg[15:0] r_54_39;
reg[15:0] r_54_40;
reg[15:0] r_54_41;
reg[15:0] r_54_42;
reg[15:0] r_54_43;
reg[15:0] r_54_44;
reg[15:0] r_54_45;
reg[15:0] r_54_46;
reg[15:0] r_54_47;
reg[15:0] r_54_48;
reg[15:0] r_54_49;
reg[15:0] r_54_50;
reg[15:0] r_54_51;
reg[15:0] r_54_52;
reg[15:0] r_54_53;
reg[15:0] r_54_54;
reg[15:0] r_54_55;
reg[15:0] r_54_56;
reg[15:0] r_54_57;
reg[15:0] r_54_58;
reg[15:0] r_54_59;
reg[15:0] r_54_60;
reg[15:0] r_54_61;
reg[15:0] r_54_62;
reg[15:0] r_54_63;
reg[15:0] r_55_0;
reg[15:0] r_55_1;
reg[15:0] r_55_2;
reg[15:0] r_55_3;
reg[15:0] r_55_4;
reg[15:0] r_55_5;
reg[15:0] r_55_6;
reg[15:0] r_55_7;
reg[15:0] r_55_8;
reg[15:0] r_55_9;
reg[15:0] r_55_10;
reg[15:0] r_55_11;
reg[15:0] r_55_12;
reg[15:0] r_55_13;
reg[15:0] r_55_14;
reg[15:0] r_55_15;
reg[15:0] r_55_16;
reg[15:0] r_55_17;
reg[15:0] r_55_18;
reg[15:0] r_55_19;
reg[15:0] r_55_20;
reg[15:0] r_55_21;
reg[15:0] r_55_22;
reg[15:0] r_55_23;
reg[15:0] r_55_24;
reg[15:0] r_55_25;
reg[15:0] r_55_26;
reg[15:0] r_55_27;
reg[15:0] r_55_28;
reg[15:0] r_55_29;
reg[15:0] r_55_30;
reg[15:0] r_55_31;
reg[15:0] r_55_32;
reg[15:0] r_55_33;
reg[15:0] r_55_34;
reg[15:0] r_55_35;
reg[15:0] r_55_36;
reg[15:0] r_55_37;
reg[15:0] r_55_38;
reg[15:0] r_55_39;
reg[15:0] r_55_40;
reg[15:0] r_55_41;
reg[15:0] r_55_42;
reg[15:0] r_55_43;
reg[15:0] r_55_44;
reg[15:0] r_55_45;
reg[15:0] r_55_46;
reg[15:0] r_55_47;
reg[15:0] r_55_48;
reg[15:0] r_55_49;
reg[15:0] r_55_50;
reg[15:0] r_55_51;
reg[15:0] r_55_52;
reg[15:0] r_55_53;
reg[15:0] r_55_54;
reg[15:0] r_55_55;
reg[15:0] r_55_56;
reg[15:0] r_55_57;
reg[15:0] r_55_58;
reg[15:0] r_55_59;
reg[15:0] r_55_60;
reg[15:0] r_55_61;
reg[15:0] r_55_62;
reg[15:0] r_55_63;
reg[15:0] r_56_0;
reg[15:0] r_56_1;
reg[15:0] r_56_2;
reg[15:0] r_56_3;
reg[15:0] r_56_4;
reg[15:0] r_56_5;
reg[15:0] r_56_6;
reg[15:0] r_56_7;
reg[15:0] r_56_8;
reg[15:0] r_56_9;
reg[15:0] r_56_10;
reg[15:0] r_56_11;
reg[15:0] r_56_12;
reg[15:0] r_56_13;
reg[15:0] r_56_14;
reg[15:0] r_56_15;
reg[15:0] r_56_16;
reg[15:0] r_56_17;
reg[15:0] r_56_18;
reg[15:0] r_56_19;
reg[15:0] r_56_20;
reg[15:0] r_56_21;
reg[15:0] r_56_22;
reg[15:0] r_56_23;
reg[15:0] r_56_24;
reg[15:0] r_56_25;
reg[15:0] r_56_26;
reg[15:0] r_56_27;
reg[15:0] r_56_28;
reg[15:0] r_56_29;
reg[15:0] r_56_30;
reg[15:0] r_56_31;
reg[15:0] r_56_32;
reg[15:0] r_56_33;
reg[15:0] r_56_34;
reg[15:0] r_56_35;
reg[15:0] r_56_36;
reg[15:0] r_56_37;
reg[15:0] r_56_38;
reg[15:0] r_56_39;
reg[15:0] r_56_40;
reg[15:0] r_56_41;
reg[15:0] r_56_42;
reg[15:0] r_56_43;
reg[15:0] r_56_44;
reg[15:0] r_56_45;
reg[15:0] r_56_46;
reg[15:0] r_56_47;
reg[15:0] r_56_48;
reg[15:0] r_56_49;
reg[15:0] r_56_50;
reg[15:0] r_56_51;
reg[15:0] r_56_52;
reg[15:0] r_56_53;
reg[15:0] r_56_54;
reg[15:0] r_56_55;
reg[15:0] r_56_56;
reg[15:0] r_56_57;
reg[15:0] r_56_58;
reg[15:0] r_56_59;
reg[15:0] r_56_60;
reg[15:0] r_56_61;
reg[15:0] r_56_62;
reg[15:0] r_56_63;
reg[15:0] r_57_0;
reg[15:0] r_57_1;
reg[15:0] r_57_2;
reg[15:0] r_57_3;
reg[15:0] r_57_4;
reg[15:0] r_57_5;
reg[15:0] r_57_6;
reg[15:0] r_57_7;
reg[15:0] r_57_8;
reg[15:0] r_57_9;
reg[15:0] r_57_10;
reg[15:0] r_57_11;
reg[15:0] r_57_12;
reg[15:0] r_57_13;
reg[15:0] r_57_14;
reg[15:0] r_57_15;
reg[15:0] r_57_16;
reg[15:0] r_57_17;
reg[15:0] r_57_18;
reg[15:0] r_57_19;
reg[15:0] r_57_20;
reg[15:0] r_57_21;
reg[15:0] r_57_22;
reg[15:0] r_57_23;
reg[15:0] r_57_24;
reg[15:0] r_57_25;
reg[15:0] r_57_26;
reg[15:0] r_57_27;
reg[15:0] r_57_28;
reg[15:0] r_57_29;
reg[15:0] r_57_30;
reg[15:0] r_57_31;
reg[15:0] r_57_32;
reg[15:0] r_57_33;
reg[15:0] r_57_34;
reg[15:0] r_57_35;
reg[15:0] r_57_36;
reg[15:0] r_57_37;
reg[15:0] r_57_38;
reg[15:0] r_57_39;
reg[15:0] r_57_40;
reg[15:0] r_57_41;
reg[15:0] r_57_42;
reg[15:0] r_57_43;
reg[15:0] r_57_44;
reg[15:0] r_57_45;
reg[15:0] r_57_46;
reg[15:0] r_57_47;
reg[15:0] r_57_48;
reg[15:0] r_57_49;
reg[15:0] r_57_50;
reg[15:0] r_57_51;
reg[15:0] r_57_52;
reg[15:0] r_57_53;
reg[15:0] r_57_54;
reg[15:0] r_57_55;
reg[15:0] r_57_56;
reg[15:0] r_57_57;
reg[15:0] r_57_58;
reg[15:0] r_57_59;
reg[15:0] r_57_60;
reg[15:0] r_57_61;
reg[15:0] r_57_62;
reg[15:0] r_57_63;
reg[15:0] r_58_0;
reg[15:0] r_58_1;
reg[15:0] r_58_2;
reg[15:0] r_58_3;
reg[15:0] r_58_4;
reg[15:0] r_58_5;
reg[15:0] r_58_6;
reg[15:0] r_58_7;
reg[15:0] r_58_8;
reg[15:0] r_58_9;
reg[15:0] r_58_10;
reg[15:0] r_58_11;
reg[15:0] r_58_12;
reg[15:0] r_58_13;
reg[15:0] r_58_14;
reg[15:0] r_58_15;
reg[15:0] r_58_16;
reg[15:0] r_58_17;
reg[15:0] r_58_18;
reg[15:0] r_58_19;
reg[15:0] r_58_20;
reg[15:0] r_58_21;
reg[15:0] r_58_22;
reg[15:0] r_58_23;
reg[15:0] r_58_24;
reg[15:0] r_58_25;
reg[15:0] r_58_26;
reg[15:0] r_58_27;
reg[15:0] r_58_28;
reg[15:0] r_58_29;
reg[15:0] r_58_30;
reg[15:0] r_58_31;
reg[15:0] r_58_32;
reg[15:0] r_58_33;
reg[15:0] r_58_34;
reg[15:0] r_58_35;
reg[15:0] r_58_36;
reg[15:0] r_58_37;
reg[15:0] r_58_38;
reg[15:0] r_58_39;
reg[15:0] r_58_40;
reg[15:0] r_58_41;
reg[15:0] r_58_42;
reg[15:0] r_58_43;
reg[15:0] r_58_44;
reg[15:0] r_58_45;
reg[15:0] r_58_46;
reg[15:0] r_58_47;
reg[15:0] r_58_48;
reg[15:0] r_58_49;
reg[15:0] r_58_50;
reg[15:0] r_58_51;
reg[15:0] r_58_52;
reg[15:0] r_58_53;
reg[15:0] r_58_54;
reg[15:0] r_58_55;
reg[15:0] r_58_56;
reg[15:0] r_58_57;
reg[15:0] r_58_58;
reg[15:0] r_58_59;
reg[15:0] r_58_60;
reg[15:0] r_58_61;
reg[15:0] r_58_62;
reg[15:0] r_58_63;
reg[15:0] r_59_0;
reg[15:0] r_59_1;
reg[15:0] r_59_2;
reg[15:0] r_59_3;
reg[15:0] r_59_4;
reg[15:0] r_59_5;
reg[15:0] r_59_6;
reg[15:0] r_59_7;
reg[15:0] r_59_8;
reg[15:0] r_59_9;
reg[15:0] r_59_10;
reg[15:0] r_59_11;
reg[15:0] r_59_12;
reg[15:0] r_59_13;
reg[15:0] r_59_14;
reg[15:0] r_59_15;
reg[15:0] r_59_16;
reg[15:0] r_59_17;
reg[15:0] r_59_18;
reg[15:0] r_59_19;
reg[15:0] r_59_20;
reg[15:0] r_59_21;
reg[15:0] r_59_22;
reg[15:0] r_59_23;
reg[15:0] r_59_24;
reg[15:0] r_59_25;
reg[15:0] r_59_26;
reg[15:0] r_59_27;
reg[15:0] r_59_28;
reg[15:0] r_59_29;
reg[15:0] r_59_30;
reg[15:0] r_59_31;
reg[15:0] r_59_32;
reg[15:0] r_59_33;
reg[15:0] r_59_34;
reg[15:0] r_59_35;
reg[15:0] r_59_36;
reg[15:0] r_59_37;
reg[15:0] r_59_38;
reg[15:0] r_59_39;
reg[15:0] r_59_40;
reg[15:0] r_59_41;
reg[15:0] r_59_42;
reg[15:0] r_59_43;
reg[15:0] r_59_44;
reg[15:0] r_59_45;
reg[15:0] r_59_46;
reg[15:0] r_59_47;
reg[15:0] r_59_48;
reg[15:0] r_59_49;
reg[15:0] r_59_50;
reg[15:0] r_59_51;
reg[15:0] r_59_52;
reg[15:0] r_59_53;
reg[15:0] r_59_54;
reg[15:0] r_59_55;
reg[15:0] r_59_56;
reg[15:0] r_59_57;
reg[15:0] r_59_58;
reg[15:0] r_59_59;
reg[15:0] r_59_60;
reg[15:0] r_59_61;
reg[15:0] r_59_62;
reg[15:0] r_59_63;
reg[15:0] r_60_0;
reg[15:0] r_60_1;
reg[15:0] r_60_2;
reg[15:0] r_60_3;
reg[15:0] r_60_4;
reg[15:0] r_60_5;
reg[15:0] r_60_6;
reg[15:0] r_60_7;
reg[15:0] r_60_8;
reg[15:0] r_60_9;
reg[15:0] r_60_10;
reg[15:0] r_60_11;
reg[15:0] r_60_12;
reg[15:0] r_60_13;
reg[15:0] r_60_14;
reg[15:0] r_60_15;
reg[15:0] r_60_16;
reg[15:0] r_60_17;
reg[15:0] r_60_18;
reg[15:0] r_60_19;
reg[15:0] r_60_20;
reg[15:0] r_60_21;
reg[15:0] r_60_22;
reg[15:0] r_60_23;
reg[15:0] r_60_24;
reg[15:0] r_60_25;
reg[15:0] r_60_26;
reg[15:0] r_60_27;
reg[15:0] r_60_28;
reg[15:0] r_60_29;
reg[15:0] r_60_30;
reg[15:0] r_60_31;
reg[15:0] r_60_32;
reg[15:0] r_60_33;
reg[15:0] r_60_34;
reg[15:0] r_60_35;
reg[15:0] r_60_36;
reg[15:0] r_60_37;
reg[15:0] r_60_38;
reg[15:0] r_60_39;
reg[15:0] r_60_40;
reg[15:0] r_60_41;
reg[15:0] r_60_42;
reg[15:0] r_60_43;
reg[15:0] r_60_44;
reg[15:0] r_60_45;
reg[15:0] r_60_46;
reg[15:0] r_60_47;
reg[15:0] r_60_48;
reg[15:0] r_60_49;
reg[15:0] r_60_50;
reg[15:0] r_60_51;
reg[15:0] r_60_52;
reg[15:0] r_60_53;
reg[15:0] r_60_54;
reg[15:0] r_60_55;
reg[15:0] r_60_56;
reg[15:0] r_60_57;
reg[15:0] r_60_58;
reg[15:0] r_60_59;
reg[15:0] r_60_60;
reg[15:0] r_60_61;
reg[15:0] r_60_62;
reg[15:0] r_60_63;
reg[15:0] r_61_0;
reg[15:0] r_61_1;
reg[15:0] r_61_2;
reg[15:0] r_61_3;
reg[15:0] r_61_4;
reg[15:0] r_61_5;
reg[15:0] r_61_6;
reg[15:0] r_61_7;
reg[15:0] r_61_8;
reg[15:0] r_61_9;
reg[15:0] r_61_10;
reg[15:0] r_61_11;
reg[15:0] r_61_12;
reg[15:0] r_61_13;
reg[15:0] r_61_14;
reg[15:0] r_61_15;
reg[15:0] r_61_16;
reg[15:0] r_61_17;
reg[15:0] r_61_18;
reg[15:0] r_61_19;
reg[15:0] r_61_20;
reg[15:0] r_61_21;
reg[15:0] r_61_22;
reg[15:0] r_61_23;
reg[15:0] r_61_24;
reg[15:0] r_61_25;
reg[15:0] r_61_26;
reg[15:0] r_61_27;
reg[15:0] r_61_28;
reg[15:0] r_61_29;
reg[15:0] r_61_30;
reg[15:0] r_61_31;
reg[15:0] r_61_32;
reg[15:0] r_61_33;
reg[15:0] r_61_34;
reg[15:0] r_61_35;
reg[15:0] r_61_36;
reg[15:0] r_61_37;
reg[15:0] r_61_38;
reg[15:0] r_61_39;
reg[15:0] r_61_40;
reg[15:0] r_61_41;
reg[15:0] r_61_42;
reg[15:0] r_61_43;
reg[15:0] r_61_44;
reg[15:0] r_61_45;
reg[15:0] r_61_46;
reg[15:0] r_61_47;
reg[15:0] r_61_48;
reg[15:0] r_61_49;
reg[15:0] r_61_50;
reg[15:0] r_61_51;
reg[15:0] r_61_52;
reg[15:0] r_61_53;
reg[15:0] r_61_54;
reg[15:0] r_61_55;
reg[15:0] r_61_56;
reg[15:0] r_61_57;
reg[15:0] r_61_58;
reg[15:0] r_61_59;
reg[15:0] r_61_60;
reg[15:0] r_61_61;
reg[15:0] r_61_62;
reg[15:0] r_61_63;
reg[15:0] r_62_0;
reg[15:0] r_62_1;
reg[15:0] r_62_2;
reg[15:0] r_62_3;
reg[15:0] r_62_4;
reg[15:0] r_62_5;
reg[15:0] r_62_6;
reg[15:0] r_62_7;
reg[15:0] r_62_8;
reg[15:0] r_62_9;
reg[15:0] r_62_10;
reg[15:0] r_62_11;
reg[15:0] r_62_12;
reg[15:0] r_62_13;
reg[15:0] r_62_14;
reg[15:0] r_62_15;
reg[15:0] r_62_16;
reg[15:0] r_62_17;
reg[15:0] r_62_18;
reg[15:0] r_62_19;
reg[15:0] r_62_20;
reg[15:0] r_62_21;
reg[15:0] r_62_22;
reg[15:0] r_62_23;
reg[15:0] r_62_24;
reg[15:0] r_62_25;
reg[15:0] r_62_26;
reg[15:0] r_62_27;
reg[15:0] r_62_28;
reg[15:0] r_62_29;
reg[15:0] r_62_30;
reg[15:0] r_62_31;
reg[15:0] r_62_32;
reg[15:0] r_62_33;
reg[15:0] r_62_34;
reg[15:0] r_62_35;
reg[15:0] r_62_36;
reg[15:0] r_62_37;
reg[15:0] r_62_38;
reg[15:0] r_62_39;
reg[15:0] r_62_40;
reg[15:0] r_62_41;
reg[15:0] r_62_42;
reg[15:0] r_62_43;
reg[15:0] r_62_44;
reg[15:0] r_62_45;
reg[15:0] r_62_46;
reg[15:0] r_62_47;
reg[15:0] r_62_48;
reg[15:0] r_62_49;
reg[15:0] r_62_50;
reg[15:0] r_62_51;
reg[15:0] r_62_52;
reg[15:0] r_62_53;
reg[15:0] r_62_54;
reg[15:0] r_62_55;
reg[15:0] r_62_56;
reg[15:0] r_62_57;
reg[15:0] r_62_58;
reg[15:0] r_62_59;
reg[15:0] r_62_60;
reg[15:0] r_62_61;
reg[15:0] r_62_62;
reg[15:0] r_62_63;
reg[15:0] r_63_0;
reg[15:0] r_63_1;
reg[15:0] r_63_2;
reg[15:0] r_63_3;
reg[15:0] r_63_4;
reg[15:0] r_63_5;
reg[15:0] r_63_6;
reg[15:0] r_63_7;
reg[15:0] r_63_8;
reg[15:0] r_63_9;
reg[15:0] r_63_10;
reg[15:0] r_63_11;
reg[15:0] r_63_12;
reg[15:0] r_63_13;
reg[15:0] r_63_14;
reg[15:0] r_63_15;
reg[15:0] r_63_16;
reg[15:0] r_63_17;
reg[15:0] r_63_18;
reg[15:0] r_63_19;
reg[15:0] r_63_20;
reg[15:0] r_63_21;
reg[15:0] r_63_22;
reg[15:0] r_63_23;
reg[15:0] r_63_24;
reg[15:0] r_63_25;
reg[15:0] r_63_26;
reg[15:0] r_63_27;
reg[15:0] r_63_28;
reg[15:0] r_63_29;
reg[15:0] r_63_30;
reg[15:0] r_63_31;
reg[15:0] r_63_32;
reg[15:0] r_63_33;
reg[15:0] r_63_34;
reg[15:0] r_63_35;
reg[15:0] r_63_36;
reg[15:0] r_63_37;
reg[15:0] r_63_38;
reg[15:0] r_63_39;
reg[15:0] r_63_40;
reg[15:0] r_63_41;
reg[15:0] r_63_42;
reg[15:0] r_63_43;
reg[15:0] r_63_44;
reg[15:0] r_63_45;
reg[15:0] r_63_46;
reg[15:0] r_63_47;
reg[15:0] r_63_48;
reg[15:0] r_63_49;
reg[15:0] r_63_50;
reg[15:0] r_63_51;
reg[15:0] r_63_52;
reg[15:0] r_63_53;
reg[15:0] r_63_54;
reg[15:0] r_63_55;
reg[15:0] r_63_56;
reg[15:0] r_63_57;
reg[15:0] r_63_58;
reg[15:0] r_63_59;
reg[15:0] r_63_60;
reg[15:0] r_63_61;
reg[15:0] r_63_62;
reg[15:0] r_63_63;
always@(posedge clk)
begin

	if (addr_selector[0]&addr_selector[0])
		data_out <= r_0_0;
		if (write_en==1'b1)
			r_0_0 <= data_in;
	if (addr_selector[0]&addr_selector[1])
		data_out <= r_0_1;
		if (write_en==1'b1)
			r_0_1 <= data_in;
	if (addr_selector[0]&addr_selector[2])
		data_out <= r_0_2;
		if (write_en==1'b1)
			r_0_2 <= data_in;
	if (addr_selector[0]&addr_selector[3])
		data_out <= r_0_3;
		if (write_en==1'b1)
			r_0_3 <= data_in;
	if (addr_selector[0]&addr_selector[4])
		data_out <= r_0_4;
		if (write_en==1'b1)
			r_0_4 <= data_in;
	if (addr_selector[0]&addr_selector[5])
		data_out <= r_0_5;
		if (write_en==1'b1)
			r_0_5 <= data_in;
	if (addr_selector[0]&addr_selector[6])
		data_out <= r_0_6;
		if (write_en==1'b1)
			r_0_6 <= data_in;
	if (addr_selector[0]&addr_selector[7])
		data_out <= r_0_7;
		if (write_en==1'b1)
			r_0_7 <= data_in;
	if (addr_selector[0]&addr_selector[8])
		data_out <= r_0_8;
		if (write_en==1'b1)
			r_0_8 <= data_in;
	if (addr_selector[0]&addr_selector[9])
		data_out <= r_0_9;
		if (write_en==1'b1)
			r_0_9 <= data_in;
	if (addr_selector[0]&addr_selector[10])
		data_out <= r_0_10;
		if (write_en==1'b1)
			r_0_10 <= data_in;
	if (addr_selector[0]&addr_selector[11])
		data_out <= r_0_11;
		if (write_en==1'b1)
			r_0_11 <= data_in;
	if (addr_selector[0]&addr_selector[12])
		data_out <= r_0_12;
		if (write_en==1'b1)
			r_0_12 <= data_in;
	if (addr_selector[0]&addr_selector[13])
		data_out <= r_0_13;
		if (write_en==1'b1)
			r_0_13 <= data_in;
	if (addr_selector[0]&addr_selector[14])
		data_out <= r_0_14;
		if (write_en==1'b1)
			r_0_14 <= data_in;
	if (addr_selector[0]&addr_selector[15])
		data_out <= r_0_15;
		if (write_en==1'b1)
			r_0_15 <= data_in;
	if (addr_selector[0]&addr_selector[16])
		data_out <= r_0_16;
		if (write_en==1'b1)
			r_0_16 <= data_in;
	if (addr_selector[0]&addr_selector[17])
		data_out <= r_0_17;
		if (write_en==1'b1)
			r_0_17 <= data_in;
	if (addr_selector[0]&addr_selector[18])
		data_out <= r_0_18;
		if (write_en==1'b1)
			r_0_18 <= data_in;
	if (addr_selector[0]&addr_selector[19])
		data_out <= r_0_19;
		if (write_en==1'b1)
			r_0_19 <= data_in;
	if (addr_selector[0]&addr_selector[20])
		data_out <= r_0_20;
		if (write_en==1'b1)
			r_0_20 <= data_in;
	if (addr_selector[0]&addr_selector[21])
		data_out <= r_0_21;
		if (write_en==1'b1)
			r_0_21 <= data_in;
	if (addr_selector[0]&addr_selector[22])
		data_out <= r_0_22;
		if (write_en==1'b1)
			r_0_22 <= data_in;
	if (addr_selector[0]&addr_selector[23])
		data_out <= r_0_23;
		if (write_en==1'b1)
			r_0_23 <= data_in;
	if (addr_selector[0]&addr_selector[24])
		data_out <= r_0_24;
		if (write_en==1'b1)
			r_0_24 <= data_in;
	if (addr_selector[0]&addr_selector[25])
		data_out <= r_0_25;
		if (write_en==1'b1)
			r_0_25 <= data_in;
	if (addr_selector[0]&addr_selector[26])
		data_out <= r_0_26;
		if (write_en==1'b1)
			r_0_26 <= data_in;
	if (addr_selector[0]&addr_selector[27])
		data_out <= r_0_27;
		if (write_en==1'b1)
			r_0_27 <= data_in;
	if (addr_selector[0]&addr_selector[28])
		data_out <= r_0_28;
		if (write_en==1'b1)
			r_0_28 <= data_in;
	if (addr_selector[0]&addr_selector[29])
		data_out <= r_0_29;
		if (write_en==1'b1)
			r_0_29 <= data_in;
	if (addr_selector[0]&addr_selector[30])
		data_out <= r_0_30;
		if (write_en==1'b1)
			r_0_30 <= data_in;
	if (addr_selector[0]&addr_selector[31])
		data_out <= r_0_31;
		if (write_en==1'b1)
			r_0_31 <= data_in;
	if (addr_selector[0]&addr_selector[32])
		data_out <= r_0_32;
		if (write_en==1'b1)
			r_0_32 <= data_in;
	if (addr_selector[0]&addr_selector[33])
		data_out <= r_0_33;
		if (write_en==1'b1)
			r_0_33 <= data_in;
	if (addr_selector[0]&addr_selector[34])
		data_out <= r_0_34;
		if (write_en==1'b1)
			r_0_34 <= data_in;
	if (addr_selector[0]&addr_selector[35])
		data_out <= r_0_35;
		if (write_en==1'b1)
			r_0_35 <= data_in;
	if (addr_selector[0]&addr_selector[36])
		data_out <= r_0_36;
		if (write_en==1'b1)
			r_0_36 <= data_in;
	if (addr_selector[0]&addr_selector[37])
		data_out <= r_0_37;
		if (write_en==1'b1)
			r_0_37 <= data_in;
	if (addr_selector[0]&addr_selector[38])
		data_out <= r_0_38;
		if (write_en==1'b1)
			r_0_38 <= data_in;
	if (addr_selector[0]&addr_selector[39])
		data_out <= r_0_39;
		if (write_en==1'b1)
			r_0_39 <= data_in;
	if (addr_selector[0]&addr_selector[40])
		data_out <= r_0_40;
		if (write_en==1'b1)
			r_0_40 <= data_in;
	if (addr_selector[0]&addr_selector[41])
		data_out <= r_0_41;
		if (write_en==1'b1)
			r_0_41 <= data_in;
	if (addr_selector[0]&addr_selector[42])
		data_out <= r_0_42;
		if (write_en==1'b1)
			r_0_42 <= data_in;
	if (addr_selector[0]&addr_selector[43])
		data_out <= r_0_43;
		if (write_en==1'b1)
			r_0_43 <= data_in;
	if (addr_selector[0]&addr_selector[44])
		data_out <= r_0_44;
		if (write_en==1'b1)
			r_0_44 <= data_in;
	if (addr_selector[0]&addr_selector[45])
		data_out <= r_0_45;
		if (write_en==1'b1)
			r_0_45 <= data_in;
	if (addr_selector[0]&addr_selector[46])
		data_out <= r_0_46;
		if (write_en==1'b1)
			r_0_46 <= data_in;
	if (addr_selector[0]&addr_selector[47])
		data_out <= r_0_47;
		if (write_en==1'b1)
			r_0_47 <= data_in;
	if (addr_selector[0]&addr_selector[48])
		data_out <= r_0_48;
		if (write_en==1'b1)
			r_0_48 <= data_in;
	if (addr_selector[0]&addr_selector[49])
		data_out <= r_0_49;
		if (write_en==1'b1)
			r_0_49 <= data_in;
	if (addr_selector[0]&addr_selector[50])
		data_out <= r_0_50;
		if (write_en==1'b1)
			r_0_50 <= data_in;
	if (addr_selector[0]&addr_selector[51])
		data_out <= r_0_51;
		if (write_en==1'b1)
			r_0_51 <= data_in;
	if (addr_selector[0]&addr_selector[52])
		data_out <= r_0_52;
		if (write_en==1'b1)
			r_0_52 <= data_in;
	if (addr_selector[0]&addr_selector[53])
		data_out <= r_0_53;
		if (write_en==1'b1)
			r_0_53 <= data_in;
	if (addr_selector[0]&addr_selector[54])
		data_out <= r_0_54;
		if (write_en==1'b1)
			r_0_54 <= data_in;
	if (addr_selector[0]&addr_selector[55])
		data_out <= r_0_55;
		if (write_en==1'b1)
			r_0_55 <= data_in;
	if (addr_selector[0]&addr_selector[56])
		data_out <= r_0_56;
		if (write_en==1'b1)
			r_0_56 <= data_in;
	if (addr_selector[0]&addr_selector[57])
		data_out <= r_0_57;
		if (write_en==1'b1)
			r_0_57 <= data_in;
	if (addr_selector[0]&addr_selector[58])
		data_out <= r_0_58;
		if (write_en==1'b1)
			r_0_58 <= data_in;
	if (addr_selector[0]&addr_selector[59])
		data_out <= r_0_59;
		if (write_en==1'b1)
			r_0_59 <= data_in;
	if (addr_selector[0]&addr_selector[60])
		data_out <= r_0_60;
		if (write_en==1'b1)
			r_0_60 <= data_in;
	if (addr_selector[0]&addr_selector[61])
		data_out <= r_0_61;
		if (write_en==1'b1)
			r_0_61 <= data_in;
	if (addr_selector[0]&addr_selector[62])
		data_out <= r_0_62;
		if (write_en==1'b1)
			r_0_62 <= data_in;
	if (addr_selector[0]&addr_selector[63])
		data_out <= r_0_63;
		if (write_en==1'b1)
			r_0_63 <= data_in;
	if (addr_selector[1]&addr_selector[0])
		data_out <= r_1_0;
		if (write_en==1'b1)
			r_1_0 <= data_in;
	if (addr_selector[1]&addr_selector[1])
		data_out <= r_1_1;
		if (write_en==1'b1)
			r_1_1 <= data_in;
	if (addr_selector[1]&addr_selector[2])
		data_out <= r_1_2;
		if (write_en==1'b1)
			r_1_2 <= data_in;
	if (addr_selector[1]&addr_selector[3])
		data_out <= r_1_3;
		if (write_en==1'b1)
			r_1_3 <= data_in;
	if (addr_selector[1]&addr_selector[4])
		data_out <= r_1_4;
		if (write_en==1'b1)
			r_1_4 <= data_in;
	if (addr_selector[1]&addr_selector[5])
		data_out <= r_1_5;
		if (write_en==1'b1)
			r_1_5 <= data_in;
	if (addr_selector[1]&addr_selector[6])
		data_out <= r_1_6;
		if (write_en==1'b1)
			r_1_6 <= data_in;
	if (addr_selector[1]&addr_selector[7])
		data_out <= r_1_7;
		if (write_en==1'b1)
			r_1_7 <= data_in;
	if (addr_selector[1]&addr_selector[8])
		data_out <= r_1_8;
		if (write_en==1'b1)
			r_1_8 <= data_in;
	if (addr_selector[1]&addr_selector[9])
		data_out <= r_1_9;
		if (write_en==1'b1)
			r_1_9 <= data_in;
	if (addr_selector[1]&addr_selector[10])
		data_out <= r_1_10;
		if (write_en==1'b1)
			r_1_10 <= data_in;
	if (addr_selector[1]&addr_selector[11])
		data_out <= r_1_11;
		if (write_en==1'b1)
			r_1_11 <= data_in;
	if (addr_selector[1]&addr_selector[12])
		data_out <= r_1_12;
		if (write_en==1'b1)
			r_1_12 <= data_in;
	if (addr_selector[1]&addr_selector[13])
		data_out <= r_1_13;
		if (write_en==1'b1)
			r_1_13 <= data_in;
	if (addr_selector[1]&addr_selector[14])
		data_out <= r_1_14;
		if (write_en==1'b1)
			r_1_14 <= data_in;
	if (addr_selector[1]&addr_selector[15])
		data_out <= r_1_15;
		if (write_en==1'b1)
			r_1_15 <= data_in;
	if (addr_selector[1]&addr_selector[16])
		data_out <= r_1_16;
		if (write_en==1'b1)
			r_1_16 <= data_in;
	if (addr_selector[1]&addr_selector[17])
		data_out <= r_1_17;
		if (write_en==1'b1)
			r_1_17 <= data_in;
	if (addr_selector[1]&addr_selector[18])
		data_out <= r_1_18;
		if (write_en==1'b1)
			r_1_18 <= data_in;
	if (addr_selector[1]&addr_selector[19])
		data_out <= r_1_19;
		if (write_en==1'b1)
			r_1_19 <= data_in;
	if (addr_selector[1]&addr_selector[20])
		data_out <= r_1_20;
		if (write_en==1'b1)
			r_1_20 <= data_in;
	if (addr_selector[1]&addr_selector[21])
		data_out <= r_1_21;
		if (write_en==1'b1)
			r_1_21 <= data_in;
	if (addr_selector[1]&addr_selector[22])
		data_out <= r_1_22;
		if (write_en==1'b1)
			r_1_22 <= data_in;
	if (addr_selector[1]&addr_selector[23])
		data_out <= r_1_23;
		if (write_en==1'b1)
			r_1_23 <= data_in;
	if (addr_selector[1]&addr_selector[24])
		data_out <= r_1_24;
		if (write_en==1'b1)
			r_1_24 <= data_in;
	if (addr_selector[1]&addr_selector[25])
		data_out <= r_1_25;
		if (write_en==1'b1)
			r_1_25 <= data_in;
	if (addr_selector[1]&addr_selector[26])
		data_out <= r_1_26;
		if (write_en==1'b1)
			r_1_26 <= data_in;
	if (addr_selector[1]&addr_selector[27])
		data_out <= r_1_27;
		if (write_en==1'b1)
			r_1_27 <= data_in;
	if (addr_selector[1]&addr_selector[28])
		data_out <= r_1_28;
		if (write_en==1'b1)
			r_1_28 <= data_in;
	if (addr_selector[1]&addr_selector[29])
		data_out <= r_1_29;
		if (write_en==1'b1)
			r_1_29 <= data_in;
	if (addr_selector[1]&addr_selector[30])
		data_out <= r_1_30;
		if (write_en==1'b1)
			r_1_30 <= data_in;
	if (addr_selector[1]&addr_selector[31])
		data_out <= r_1_31;
		if (write_en==1'b1)
			r_1_31 <= data_in;
	if (addr_selector[1]&addr_selector[32])
		data_out <= r_1_32;
		if (write_en==1'b1)
			r_1_32 <= data_in;
	if (addr_selector[1]&addr_selector[33])
		data_out <= r_1_33;
		if (write_en==1'b1)
			r_1_33 <= data_in;
	if (addr_selector[1]&addr_selector[34])
		data_out <= r_1_34;
		if (write_en==1'b1)
			r_1_34 <= data_in;
	if (addr_selector[1]&addr_selector[35])
		data_out <= r_1_35;
		if (write_en==1'b1)
			r_1_35 <= data_in;
	if (addr_selector[1]&addr_selector[36])
		data_out <= r_1_36;
		if (write_en==1'b1)
			r_1_36 <= data_in;
	if (addr_selector[1]&addr_selector[37])
		data_out <= r_1_37;
		if (write_en==1'b1)
			r_1_37 <= data_in;
	if (addr_selector[1]&addr_selector[38])
		data_out <= r_1_38;
		if (write_en==1'b1)
			r_1_38 <= data_in;
	if (addr_selector[1]&addr_selector[39])
		data_out <= r_1_39;
		if (write_en==1'b1)
			r_1_39 <= data_in;
	if (addr_selector[1]&addr_selector[40])
		data_out <= r_1_40;
		if (write_en==1'b1)
			r_1_40 <= data_in;
	if (addr_selector[1]&addr_selector[41])
		data_out <= r_1_41;
		if (write_en==1'b1)
			r_1_41 <= data_in;
	if (addr_selector[1]&addr_selector[42])
		data_out <= r_1_42;
		if (write_en==1'b1)
			r_1_42 <= data_in;
	if (addr_selector[1]&addr_selector[43])
		data_out <= r_1_43;
		if (write_en==1'b1)
			r_1_43 <= data_in;
	if (addr_selector[1]&addr_selector[44])
		data_out <= r_1_44;
		if (write_en==1'b1)
			r_1_44 <= data_in;
	if (addr_selector[1]&addr_selector[45])
		data_out <= r_1_45;
		if (write_en==1'b1)
			r_1_45 <= data_in;
	if (addr_selector[1]&addr_selector[46])
		data_out <= r_1_46;
		if (write_en==1'b1)
			r_1_46 <= data_in;
	if (addr_selector[1]&addr_selector[47])
		data_out <= r_1_47;
		if (write_en==1'b1)
			r_1_47 <= data_in;
	if (addr_selector[1]&addr_selector[48])
		data_out <= r_1_48;
		if (write_en==1'b1)
			r_1_48 <= data_in;
	if (addr_selector[1]&addr_selector[49])
		data_out <= r_1_49;
		if (write_en==1'b1)
			r_1_49 <= data_in;
	if (addr_selector[1]&addr_selector[50])
		data_out <= r_1_50;
		if (write_en==1'b1)
			r_1_50 <= data_in;
	if (addr_selector[1]&addr_selector[51])
		data_out <= r_1_51;
		if (write_en==1'b1)
			r_1_51 <= data_in;
	if (addr_selector[1]&addr_selector[52])
		data_out <= r_1_52;
		if (write_en==1'b1)
			r_1_52 <= data_in;
	if (addr_selector[1]&addr_selector[53])
		data_out <= r_1_53;
		if (write_en==1'b1)
			r_1_53 <= data_in;
	if (addr_selector[1]&addr_selector[54])
		data_out <= r_1_54;
		if (write_en==1'b1)
			r_1_54 <= data_in;
	if (addr_selector[1]&addr_selector[55])
		data_out <= r_1_55;
		if (write_en==1'b1)
			r_1_55 <= data_in;
	if (addr_selector[1]&addr_selector[56])
		data_out <= r_1_56;
		if (write_en==1'b1)
			r_1_56 <= data_in;
	if (addr_selector[1]&addr_selector[57])
		data_out <= r_1_57;
		if (write_en==1'b1)
			r_1_57 <= data_in;
	if (addr_selector[1]&addr_selector[58])
		data_out <= r_1_58;
		if (write_en==1'b1)
			r_1_58 <= data_in;
	if (addr_selector[1]&addr_selector[59])
		data_out <= r_1_59;
		if (write_en==1'b1)
			r_1_59 <= data_in;
	if (addr_selector[1]&addr_selector[60])
		data_out <= r_1_60;
		if (write_en==1'b1)
			r_1_60 <= data_in;
	if (addr_selector[1]&addr_selector[61])
		data_out <= r_1_61;
		if (write_en==1'b1)
			r_1_61 <= data_in;
	if (addr_selector[1]&addr_selector[62])
		data_out <= r_1_62;
		if (write_en==1'b1)
			r_1_62 <= data_in;
	if (addr_selector[1]&addr_selector[63])
		data_out <= r_1_63;
		if (write_en==1'b1)
			r_1_63 <= data_in;
	if (addr_selector[2]&addr_selector[0])
		data_out <= r_2_0;
		if (write_en==1'b1)
			r_2_0 <= data_in;
	if (addr_selector[2]&addr_selector[1])
		data_out <= r_2_1;
		if (write_en==1'b1)
			r_2_1 <= data_in;
	if (addr_selector[2]&addr_selector[2])
		data_out <= r_2_2;
		if (write_en==1'b1)
			r_2_2 <= data_in;
	if (addr_selector[2]&addr_selector[3])
		data_out <= r_2_3;
		if (write_en==1'b1)
			r_2_3 <= data_in;
	if (addr_selector[2]&addr_selector[4])
		data_out <= r_2_4;
		if (write_en==1'b1)
			r_2_4 <= data_in;
	if (addr_selector[2]&addr_selector[5])
		data_out <= r_2_5;
		if (write_en==1'b1)
			r_2_5 <= data_in;
	if (addr_selector[2]&addr_selector[6])
		data_out <= r_2_6;
		if (write_en==1'b1)
			r_2_6 <= data_in;
	if (addr_selector[2]&addr_selector[7])
		data_out <= r_2_7;
		if (write_en==1'b1)
			r_2_7 <= data_in;
	if (addr_selector[2]&addr_selector[8])
		data_out <= r_2_8;
		if (write_en==1'b1)
			r_2_8 <= data_in;
	if (addr_selector[2]&addr_selector[9])
		data_out <= r_2_9;
		if (write_en==1'b1)
			r_2_9 <= data_in;
	if (addr_selector[2]&addr_selector[10])
		data_out <= r_2_10;
		if (write_en==1'b1)
			r_2_10 <= data_in;
	if (addr_selector[2]&addr_selector[11])
		data_out <= r_2_11;
		if (write_en==1'b1)
			r_2_11 <= data_in;
	if (addr_selector[2]&addr_selector[12])
		data_out <= r_2_12;
		if (write_en==1'b1)
			r_2_12 <= data_in;
	if (addr_selector[2]&addr_selector[13])
		data_out <= r_2_13;
		if (write_en==1'b1)
			r_2_13 <= data_in;
	if (addr_selector[2]&addr_selector[14])
		data_out <= r_2_14;
		if (write_en==1'b1)
			r_2_14 <= data_in;
	if (addr_selector[2]&addr_selector[15])
		data_out <= r_2_15;
		if (write_en==1'b1)
			r_2_15 <= data_in;
	if (addr_selector[2]&addr_selector[16])
		data_out <= r_2_16;
		if (write_en==1'b1)
			r_2_16 <= data_in;
	if (addr_selector[2]&addr_selector[17])
		data_out <= r_2_17;
		if (write_en==1'b1)
			r_2_17 <= data_in;
	if (addr_selector[2]&addr_selector[18])
		data_out <= r_2_18;
		if (write_en==1'b1)
			r_2_18 <= data_in;
	if (addr_selector[2]&addr_selector[19])
		data_out <= r_2_19;
		if (write_en==1'b1)
			r_2_19 <= data_in;
	if (addr_selector[2]&addr_selector[20])
		data_out <= r_2_20;
		if (write_en==1'b1)
			r_2_20 <= data_in;
	if (addr_selector[2]&addr_selector[21])
		data_out <= r_2_21;
		if (write_en==1'b1)
			r_2_21 <= data_in;
	if (addr_selector[2]&addr_selector[22])
		data_out <= r_2_22;
		if (write_en==1'b1)
			r_2_22 <= data_in;
	if (addr_selector[2]&addr_selector[23])
		data_out <= r_2_23;
		if (write_en==1'b1)
			r_2_23 <= data_in;
	if (addr_selector[2]&addr_selector[24])
		data_out <= r_2_24;
		if (write_en==1'b1)
			r_2_24 <= data_in;
	if (addr_selector[2]&addr_selector[25])
		data_out <= r_2_25;
		if (write_en==1'b1)
			r_2_25 <= data_in;
	if (addr_selector[2]&addr_selector[26])
		data_out <= r_2_26;
		if (write_en==1'b1)
			r_2_26 <= data_in;
	if (addr_selector[2]&addr_selector[27])
		data_out <= r_2_27;
		if (write_en==1'b1)
			r_2_27 <= data_in;
	if (addr_selector[2]&addr_selector[28])
		data_out <= r_2_28;
		if (write_en==1'b1)
			r_2_28 <= data_in;
	if (addr_selector[2]&addr_selector[29])
		data_out <= r_2_29;
		if (write_en==1'b1)
			r_2_29 <= data_in;
	if (addr_selector[2]&addr_selector[30])
		data_out <= r_2_30;
		if (write_en==1'b1)
			r_2_30 <= data_in;
	if (addr_selector[2]&addr_selector[31])
		data_out <= r_2_31;
		if (write_en==1'b1)
			r_2_31 <= data_in;
	if (addr_selector[2]&addr_selector[32])
		data_out <= r_2_32;
		if (write_en==1'b1)
			r_2_32 <= data_in;
	if (addr_selector[2]&addr_selector[33])
		data_out <= r_2_33;
		if (write_en==1'b1)
			r_2_33 <= data_in;
	if (addr_selector[2]&addr_selector[34])
		data_out <= r_2_34;
		if (write_en==1'b1)
			r_2_34 <= data_in;
	if (addr_selector[2]&addr_selector[35])
		data_out <= r_2_35;
		if (write_en==1'b1)
			r_2_35 <= data_in;
	if (addr_selector[2]&addr_selector[36])
		data_out <= r_2_36;
		if (write_en==1'b1)
			r_2_36 <= data_in;
	if (addr_selector[2]&addr_selector[37])
		data_out <= r_2_37;
		if (write_en==1'b1)
			r_2_37 <= data_in;
	if (addr_selector[2]&addr_selector[38])
		data_out <= r_2_38;
		if (write_en==1'b1)
			r_2_38 <= data_in;
	if (addr_selector[2]&addr_selector[39])
		data_out <= r_2_39;
		if (write_en==1'b1)
			r_2_39 <= data_in;
	if (addr_selector[2]&addr_selector[40])
		data_out <= r_2_40;
		if (write_en==1'b1)
			r_2_40 <= data_in;
	if (addr_selector[2]&addr_selector[41])
		data_out <= r_2_41;
		if (write_en==1'b1)
			r_2_41 <= data_in;
	if (addr_selector[2]&addr_selector[42])
		data_out <= r_2_42;
		if (write_en==1'b1)
			r_2_42 <= data_in;
	if (addr_selector[2]&addr_selector[43])
		data_out <= r_2_43;
		if (write_en==1'b1)
			r_2_43 <= data_in;
	if (addr_selector[2]&addr_selector[44])
		data_out <= r_2_44;
		if (write_en==1'b1)
			r_2_44 <= data_in;
	if (addr_selector[2]&addr_selector[45])
		data_out <= r_2_45;
		if (write_en==1'b1)
			r_2_45 <= data_in;
	if (addr_selector[2]&addr_selector[46])
		data_out <= r_2_46;
		if (write_en==1'b1)
			r_2_46 <= data_in;
	if (addr_selector[2]&addr_selector[47])
		data_out <= r_2_47;
		if (write_en==1'b1)
			r_2_47 <= data_in;
	if (addr_selector[2]&addr_selector[48])
		data_out <= r_2_48;
		if (write_en==1'b1)
			r_2_48 <= data_in;
	if (addr_selector[2]&addr_selector[49])
		data_out <= r_2_49;
		if (write_en==1'b1)
			r_2_49 <= data_in;
	if (addr_selector[2]&addr_selector[50])
		data_out <= r_2_50;
		if (write_en==1'b1)
			r_2_50 <= data_in;
	if (addr_selector[2]&addr_selector[51])
		data_out <= r_2_51;
		if (write_en==1'b1)
			r_2_51 <= data_in;
	if (addr_selector[2]&addr_selector[52])
		data_out <= r_2_52;
		if (write_en==1'b1)
			r_2_52 <= data_in;
	if (addr_selector[2]&addr_selector[53])
		data_out <= r_2_53;
		if (write_en==1'b1)
			r_2_53 <= data_in;
	if (addr_selector[2]&addr_selector[54])
		data_out <= r_2_54;
		if (write_en==1'b1)
			r_2_54 <= data_in;
	if (addr_selector[2]&addr_selector[55])
		data_out <= r_2_55;
		if (write_en==1'b1)
			r_2_55 <= data_in;
	if (addr_selector[2]&addr_selector[56])
		data_out <= r_2_56;
		if (write_en==1'b1)
			r_2_56 <= data_in;
	if (addr_selector[2]&addr_selector[57])
		data_out <= r_2_57;
		if (write_en==1'b1)
			r_2_57 <= data_in;
	if (addr_selector[2]&addr_selector[58])
		data_out <= r_2_58;
		if (write_en==1'b1)
			r_2_58 <= data_in;
	if (addr_selector[2]&addr_selector[59])
		data_out <= r_2_59;
		if (write_en==1'b1)
			r_2_59 <= data_in;
	if (addr_selector[2]&addr_selector[60])
		data_out <= r_2_60;
		if (write_en==1'b1)
			r_2_60 <= data_in;
	if (addr_selector[2]&addr_selector[61])
		data_out <= r_2_61;
		if (write_en==1'b1)
			r_2_61 <= data_in;
	if (addr_selector[2]&addr_selector[62])
		data_out <= r_2_62;
		if (write_en==1'b1)
			r_2_62 <= data_in;
	if (addr_selector[2]&addr_selector[63])
		data_out <= r_2_63;
		if (write_en==1'b1)
			r_2_63 <= data_in;
	if (addr_selector[3]&addr_selector[0])
		data_out <= r_3_0;
		if (write_en==1'b1)
			r_3_0 <= data_in;
	if (addr_selector[3]&addr_selector[1])
		data_out <= r_3_1;
		if (write_en==1'b1)
			r_3_1 <= data_in;
	if (addr_selector[3]&addr_selector[2])
		data_out <= r_3_2;
		if (write_en==1'b1)
			r_3_2 <= data_in;
	if (addr_selector[3]&addr_selector[3])
		data_out <= r_3_3;
		if (write_en==1'b1)
			r_3_3 <= data_in;
	if (addr_selector[3]&addr_selector[4])
		data_out <= r_3_4;
		if (write_en==1'b1)
			r_3_4 <= data_in;
	if (addr_selector[3]&addr_selector[5])
		data_out <= r_3_5;
		if (write_en==1'b1)
			r_3_5 <= data_in;
	if (addr_selector[3]&addr_selector[6])
		data_out <= r_3_6;
		if (write_en==1'b1)
			r_3_6 <= data_in;
	if (addr_selector[3]&addr_selector[7])
		data_out <= r_3_7;
		if (write_en==1'b1)
			r_3_7 <= data_in;
	if (addr_selector[3]&addr_selector[8])
		data_out <= r_3_8;
		if (write_en==1'b1)
			r_3_8 <= data_in;
	if (addr_selector[3]&addr_selector[9])
		data_out <= r_3_9;
		if (write_en==1'b1)
			r_3_9 <= data_in;
	if (addr_selector[3]&addr_selector[10])
		data_out <= r_3_10;
		if (write_en==1'b1)
			r_3_10 <= data_in;
	if (addr_selector[3]&addr_selector[11])
		data_out <= r_3_11;
		if (write_en==1'b1)
			r_3_11 <= data_in;
	if (addr_selector[3]&addr_selector[12])
		data_out <= r_3_12;
		if (write_en==1'b1)
			r_3_12 <= data_in;
	if (addr_selector[3]&addr_selector[13])
		data_out <= r_3_13;
		if (write_en==1'b1)
			r_3_13 <= data_in;
	if (addr_selector[3]&addr_selector[14])
		data_out <= r_3_14;
		if (write_en==1'b1)
			r_3_14 <= data_in;
	if (addr_selector[3]&addr_selector[15])
		data_out <= r_3_15;
		if (write_en==1'b1)
			r_3_15 <= data_in;
	if (addr_selector[3]&addr_selector[16])
		data_out <= r_3_16;
		if (write_en==1'b1)
			r_3_16 <= data_in;
	if (addr_selector[3]&addr_selector[17])
		data_out <= r_3_17;
		if (write_en==1'b1)
			r_3_17 <= data_in;
	if (addr_selector[3]&addr_selector[18])
		data_out <= r_3_18;
		if (write_en==1'b1)
			r_3_18 <= data_in;
	if (addr_selector[3]&addr_selector[19])
		data_out <= r_3_19;
		if (write_en==1'b1)
			r_3_19 <= data_in;
	if (addr_selector[3]&addr_selector[20])
		data_out <= r_3_20;
		if (write_en==1'b1)
			r_3_20 <= data_in;
	if (addr_selector[3]&addr_selector[21])
		data_out <= r_3_21;
		if (write_en==1'b1)
			r_3_21 <= data_in;
	if (addr_selector[3]&addr_selector[22])
		data_out <= r_3_22;
		if (write_en==1'b1)
			r_3_22 <= data_in;
	if (addr_selector[3]&addr_selector[23])
		data_out <= r_3_23;
		if (write_en==1'b1)
			r_3_23 <= data_in;
	if (addr_selector[3]&addr_selector[24])
		data_out <= r_3_24;
		if (write_en==1'b1)
			r_3_24 <= data_in;
	if (addr_selector[3]&addr_selector[25])
		data_out <= r_3_25;
		if (write_en==1'b1)
			r_3_25 <= data_in;
	if (addr_selector[3]&addr_selector[26])
		data_out <= r_3_26;
		if (write_en==1'b1)
			r_3_26 <= data_in;
	if (addr_selector[3]&addr_selector[27])
		data_out <= r_3_27;
		if (write_en==1'b1)
			r_3_27 <= data_in;
	if (addr_selector[3]&addr_selector[28])
		data_out <= r_3_28;
		if (write_en==1'b1)
			r_3_28 <= data_in;
	if (addr_selector[3]&addr_selector[29])
		data_out <= r_3_29;
		if (write_en==1'b1)
			r_3_29 <= data_in;
	if (addr_selector[3]&addr_selector[30])
		data_out <= r_3_30;
		if (write_en==1'b1)
			r_3_30 <= data_in;
	if (addr_selector[3]&addr_selector[31])
		data_out <= r_3_31;
		if (write_en==1'b1)
			r_3_31 <= data_in;
	if (addr_selector[3]&addr_selector[32])
		data_out <= r_3_32;
		if (write_en==1'b1)
			r_3_32 <= data_in;
	if (addr_selector[3]&addr_selector[33])
		data_out <= r_3_33;
		if (write_en==1'b1)
			r_3_33 <= data_in;
	if (addr_selector[3]&addr_selector[34])
		data_out <= r_3_34;
		if (write_en==1'b1)
			r_3_34 <= data_in;
	if (addr_selector[3]&addr_selector[35])
		data_out <= r_3_35;
		if (write_en==1'b1)
			r_3_35 <= data_in;
	if (addr_selector[3]&addr_selector[36])
		data_out <= r_3_36;
		if (write_en==1'b1)
			r_3_36 <= data_in;
	if (addr_selector[3]&addr_selector[37])
		data_out <= r_3_37;
		if (write_en==1'b1)
			r_3_37 <= data_in;
	if (addr_selector[3]&addr_selector[38])
		data_out <= r_3_38;
		if (write_en==1'b1)
			r_3_38 <= data_in;
	if (addr_selector[3]&addr_selector[39])
		data_out <= r_3_39;
		if (write_en==1'b1)
			r_3_39 <= data_in;
	if (addr_selector[3]&addr_selector[40])
		data_out <= r_3_40;
		if (write_en==1'b1)
			r_3_40 <= data_in;
	if (addr_selector[3]&addr_selector[41])
		data_out <= r_3_41;
		if (write_en==1'b1)
			r_3_41 <= data_in;
	if (addr_selector[3]&addr_selector[42])
		data_out <= r_3_42;
		if (write_en==1'b1)
			r_3_42 <= data_in;
	if (addr_selector[3]&addr_selector[43])
		data_out <= r_3_43;
		if (write_en==1'b1)
			r_3_43 <= data_in;
	if (addr_selector[3]&addr_selector[44])
		data_out <= r_3_44;
		if (write_en==1'b1)
			r_3_44 <= data_in;
	if (addr_selector[3]&addr_selector[45])
		data_out <= r_3_45;
		if (write_en==1'b1)
			r_3_45 <= data_in;
	if (addr_selector[3]&addr_selector[46])
		data_out <= r_3_46;
		if (write_en==1'b1)
			r_3_46 <= data_in;
	if (addr_selector[3]&addr_selector[47])
		data_out <= r_3_47;
		if (write_en==1'b1)
			r_3_47 <= data_in;
	if (addr_selector[3]&addr_selector[48])
		data_out <= r_3_48;
		if (write_en==1'b1)
			r_3_48 <= data_in;
	if (addr_selector[3]&addr_selector[49])
		data_out <= r_3_49;
		if (write_en==1'b1)
			r_3_49 <= data_in;
	if (addr_selector[3]&addr_selector[50])
		data_out <= r_3_50;
		if (write_en==1'b1)
			r_3_50 <= data_in;
	if (addr_selector[3]&addr_selector[51])
		data_out <= r_3_51;
		if (write_en==1'b1)
			r_3_51 <= data_in;
	if (addr_selector[3]&addr_selector[52])
		data_out <= r_3_52;
		if (write_en==1'b1)
			r_3_52 <= data_in;
	if (addr_selector[3]&addr_selector[53])
		data_out <= r_3_53;
		if (write_en==1'b1)
			r_3_53 <= data_in;
	if (addr_selector[3]&addr_selector[54])
		data_out <= r_3_54;
		if (write_en==1'b1)
			r_3_54 <= data_in;
	if (addr_selector[3]&addr_selector[55])
		data_out <= r_3_55;
		if (write_en==1'b1)
			r_3_55 <= data_in;
	if (addr_selector[3]&addr_selector[56])
		data_out <= r_3_56;
		if (write_en==1'b1)
			r_3_56 <= data_in;
	if (addr_selector[3]&addr_selector[57])
		data_out <= r_3_57;
		if (write_en==1'b1)
			r_3_57 <= data_in;
	if (addr_selector[3]&addr_selector[58])
		data_out <= r_3_58;
		if (write_en==1'b1)
			r_3_58 <= data_in;
	if (addr_selector[3]&addr_selector[59])
		data_out <= r_3_59;
		if (write_en==1'b1)
			r_3_59 <= data_in;
	if (addr_selector[3]&addr_selector[60])
		data_out <= r_3_60;
		if (write_en==1'b1)
			r_3_60 <= data_in;
	if (addr_selector[3]&addr_selector[61])
		data_out <= r_3_61;
		if (write_en==1'b1)
			r_3_61 <= data_in;
	if (addr_selector[3]&addr_selector[62])
		data_out <= r_3_62;
		if (write_en==1'b1)
			r_3_62 <= data_in;
	if (addr_selector[3]&addr_selector[63])
		data_out <= r_3_63;
		if (write_en==1'b1)
			r_3_63 <= data_in;
	if (addr_selector[4]&addr_selector[0])
		data_out <= r_4_0;
		if (write_en==1'b1)
			r_4_0 <= data_in;
	if (addr_selector[4]&addr_selector[1])
		data_out <= r_4_1;
		if (write_en==1'b1)
			r_4_1 <= data_in;
	if (addr_selector[4]&addr_selector[2])
		data_out <= r_4_2;
		if (write_en==1'b1)
			r_4_2 <= data_in;
	if (addr_selector[4]&addr_selector[3])
		data_out <= r_4_3;
		if (write_en==1'b1)
			r_4_3 <= data_in;
	if (addr_selector[4]&addr_selector[4])
		data_out <= r_4_4;
		if (write_en==1'b1)
			r_4_4 <= data_in;
	if (addr_selector[4]&addr_selector[5])
		data_out <= r_4_5;
		if (write_en==1'b1)
			r_4_5 <= data_in;
	if (addr_selector[4]&addr_selector[6])
		data_out <= r_4_6;
		if (write_en==1'b1)
			r_4_6 <= data_in;
	if (addr_selector[4]&addr_selector[7])
		data_out <= r_4_7;
		if (write_en==1'b1)
			r_4_7 <= data_in;
	if (addr_selector[4]&addr_selector[8])
		data_out <= r_4_8;
		if (write_en==1'b1)
			r_4_8 <= data_in;
	if (addr_selector[4]&addr_selector[9])
		data_out <= r_4_9;
		if (write_en==1'b1)
			r_4_9 <= data_in;
	if (addr_selector[4]&addr_selector[10])
		data_out <= r_4_10;
		if (write_en==1'b1)
			r_4_10 <= data_in;
	if (addr_selector[4]&addr_selector[11])
		data_out <= r_4_11;
		if (write_en==1'b1)
			r_4_11 <= data_in;
	if (addr_selector[4]&addr_selector[12])
		data_out <= r_4_12;
		if (write_en==1'b1)
			r_4_12 <= data_in;
	if (addr_selector[4]&addr_selector[13])
		data_out <= r_4_13;
		if (write_en==1'b1)
			r_4_13 <= data_in;
	if (addr_selector[4]&addr_selector[14])
		data_out <= r_4_14;
		if (write_en==1'b1)
			r_4_14 <= data_in;
	if (addr_selector[4]&addr_selector[15])
		data_out <= r_4_15;
		if (write_en==1'b1)
			r_4_15 <= data_in;
	if (addr_selector[4]&addr_selector[16])
		data_out <= r_4_16;
		if (write_en==1'b1)
			r_4_16 <= data_in;
	if (addr_selector[4]&addr_selector[17])
		data_out <= r_4_17;
		if (write_en==1'b1)
			r_4_17 <= data_in;
	if (addr_selector[4]&addr_selector[18])
		data_out <= r_4_18;
		if (write_en==1'b1)
			r_4_18 <= data_in;
	if (addr_selector[4]&addr_selector[19])
		data_out <= r_4_19;
		if (write_en==1'b1)
			r_4_19 <= data_in;
	if (addr_selector[4]&addr_selector[20])
		data_out <= r_4_20;
		if (write_en==1'b1)
			r_4_20 <= data_in;
	if (addr_selector[4]&addr_selector[21])
		data_out <= r_4_21;
		if (write_en==1'b1)
			r_4_21 <= data_in;
	if (addr_selector[4]&addr_selector[22])
		data_out <= r_4_22;
		if (write_en==1'b1)
			r_4_22 <= data_in;
	if (addr_selector[4]&addr_selector[23])
		data_out <= r_4_23;
		if (write_en==1'b1)
			r_4_23 <= data_in;
	if (addr_selector[4]&addr_selector[24])
		data_out <= r_4_24;
		if (write_en==1'b1)
			r_4_24 <= data_in;
	if (addr_selector[4]&addr_selector[25])
		data_out <= r_4_25;
		if (write_en==1'b1)
			r_4_25 <= data_in;
	if (addr_selector[4]&addr_selector[26])
		data_out <= r_4_26;
		if (write_en==1'b1)
			r_4_26 <= data_in;
	if (addr_selector[4]&addr_selector[27])
		data_out <= r_4_27;
		if (write_en==1'b1)
			r_4_27 <= data_in;
	if (addr_selector[4]&addr_selector[28])
		data_out <= r_4_28;
		if (write_en==1'b1)
			r_4_28 <= data_in;
	if (addr_selector[4]&addr_selector[29])
		data_out <= r_4_29;
		if (write_en==1'b1)
			r_4_29 <= data_in;
	if (addr_selector[4]&addr_selector[30])
		data_out <= r_4_30;
		if (write_en==1'b1)
			r_4_30 <= data_in;
	if (addr_selector[4]&addr_selector[31])
		data_out <= r_4_31;
		if (write_en==1'b1)
			r_4_31 <= data_in;
	if (addr_selector[4]&addr_selector[32])
		data_out <= r_4_32;
		if (write_en==1'b1)
			r_4_32 <= data_in;
	if (addr_selector[4]&addr_selector[33])
		data_out <= r_4_33;
		if (write_en==1'b1)
			r_4_33 <= data_in;
	if (addr_selector[4]&addr_selector[34])
		data_out <= r_4_34;
		if (write_en==1'b1)
			r_4_34 <= data_in;
	if (addr_selector[4]&addr_selector[35])
		data_out <= r_4_35;
		if (write_en==1'b1)
			r_4_35 <= data_in;
	if (addr_selector[4]&addr_selector[36])
		data_out <= r_4_36;
		if (write_en==1'b1)
			r_4_36 <= data_in;
	if (addr_selector[4]&addr_selector[37])
		data_out <= r_4_37;
		if (write_en==1'b1)
			r_4_37 <= data_in;
	if (addr_selector[4]&addr_selector[38])
		data_out <= r_4_38;
		if (write_en==1'b1)
			r_4_38 <= data_in;
	if (addr_selector[4]&addr_selector[39])
		data_out <= r_4_39;
		if (write_en==1'b1)
			r_4_39 <= data_in;
	if (addr_selector[4]&addr_selector[40])
		data_out <= r_4_40;
		if (write_en==1'b1)
			r_4_40 <= data_in;
	if (addr_selector[4]&addr_selector[41])
		data_out <= r_4_41;
		if (write_en==1'b1)
			r_4_41 <= data_in;
	if (addr_selector[4]&addr_selector[42])
		data_out <= r_4_42;
		if (write_en==1'b1)
			r_4_42 <= data_in;
	if (addr_selector[4]&addr_selector[43])
		data_out <= r_4_43;
		if (write_en==1'b1)
			r_4_43 <= data_in;
	if (addr_selector[4]&addr_selector[44])
		data_out <= r_4_44;
		if (write_en==1'b1)
			r_4_44 <= data_in;
	if (addr_selector[4]&addr_selector[45])
		data_out <= r_4_45;
		if (write_en==1'b1)
			r_4_45 <= data_in;
	if (addr_selector[4]&addr_selector[46])
		data_out <= r_4_46;
		if (write_en==1'b1)
			r_4_46 <= data_in;
	if (addr_selector[4]&addr_selector[47])
		data_out <= r_4_47;
		if (write_en==1'b1)
			r_4_47 <= data_in;
	if (addr_selector[4]&addr_selector[48])
		data_out <= r_4_48;
		if (write_en==1'b1)
			r_4_48 <= data_in;
	if (addr_selector[4]&addr_selector[49])
		data_out <= r_4_49;
		if (write_en==1'b1)
			r_4_49 <= data_in;
	if (addr_selector[4]&addr_selector[50])
		data_out <= r_4_50;
		if (write_en==1'b1)
			r_4_50 <= data_in;
	if (addr_selector[4]&addr_selector[51])
		data_out <= r_4_51;
		if (write_en==1'b1)
			r_4_51 <= data_in;
	if (addr_selector[4]&addr_selector[52])
		data_out <= r_4_52;
		if (write_en==1'b1)
			r_4_52 <= data_in;
	if (addr_selector[4]&addr_selector[53])
		data_out <= r_4_53;
		if (write_en==1'b1)
			r_4_53 <= data_in;
	if (addr_selector[4]&addr_selector[54])
		data_out <= r_4_54;
		if (write_en==1'b1)
			r_4_54 <= data_in;
	if (addr_selector[4]&addr_selector[55])
		data_out <= r_4_55;
		if (write_en==1'b1)
			r_4_55 <= data_in;
	if (addr_selector[4]&addr_selector[56])
		data_out <= r_4_56;
		if (write_en==1'b1)
			r_4_56 <= data_in;
	if (addr_selector[4]&addr_selector[57])
		data_out <= r_4_57;
		if (write_en==1'b1)
			r_4_57 <= data_in;
	if (addr_selector[4]&addr_selector[58])
		data_out <= r_4_58;
		if (write_en==1'b1)
			r_4_58 <= data_in;
	if (addr_selector[4]&addr_selector[59])
		data_out <= r_4_59;
		if (write_en==1'b1)
			r_4_59 <= data_in;
	if (addr_selector[4]&addr_selector[60])
		data_out <= r_4_60;
		if (write_en==1'b1)
			r_4_60 <= data_in;
	if (addr_selector[4]&addr_selector[61])
		data_out <= r_4_61;
		if (write_en==1'b1)
			r_4_61 <= data_in;
	if (addr_selector[4]&addr_selector[62])
		data_out <= r_4_62;
		if (write_en==1'b1)
			r_4_62 <= data_in;
	if (addr_selector[4]&addr_selector[63])
		data_out <= r_4_63;
		if (write_en==1'b1)
			r_4_63 <= data_in;
	if (addr_selector[5]&addr_selector[0])
		data_out <= r_5_0;
		if (write_en==1'b1)
			r_5_0 <= data_in;
	if (addr_selector[5]&addr_selector[1])
		data_out <= r_5_1;
		if (write_en==1'b1)
			r_5_1 <= data_in;
	if (addr_selector[5]&addr_selector[2])
		data_out <= r_5_2;
		if (write_en==1'b1)
			r_5_2 <= data_in;
	if (addr_selector[5]&addr_selector[3])
		data_out <= r_5_3;
		if (write_en==1'b1)
			r_5_3 <= data_in;
	if (addr_selector[5]&addr_selector[4])
		data_out <= r_5_4;
		if (write_en==1'b1)
			r_5_4 <= data_in;
	if (addr_selector[5]&addr_selector[5])
		data_out <= r_5_5;
		if (write_en==1'b1)
			r_5_5 <= data_in;
	if (addr_selector[5]&addr_selector[6])
		data_out <= r_5_6;
		if (write_en==1'b1)
			r_5_6 <= data_in;
	if (addr_selector[5]&addr_selector[7])
		data_out <= r_5_7;
		if (write_en==1'b1)
			r_5_7 <= data_in;
	if (addr_selector[5]&addr_selector[8])
		data_out <= r_5_8;
		if (write_en==1'b1)
			r_5_8 <= data_in;
	if (addr_selector[5]&addr_selector[9])
		data_out <= r_5_9;
		if (write_en==1'b1)
			r_5_9 <= data_in;
	if (addr_selector[5]&addr_selector[10])
		data_out <= r_5_10;
		if (write_en==1'b1)
			r_5_10 <= data_in;
	if (addr_selector[5]&addr_selector[11])
		data_out <= r_5_11;
		if (write_en==1'b1)
			r_5_11 <= data_in;
	if (addr_selector[5]&addr_selector[12])
		data_out <= r_5_12;
		if (write_en==1'b1)
			r_5_12 <= data_in;
	if (addr_selector[5]&addr_selector[13])
		data_out <= r_5_13;
		if (write_en==1'b1)
			r_5_13 <= data_in;
	if (addr_selector[5]&addr_selector[14])
		data_out <= r_5_14;
		if (write_en==1'b1)
			r_5_14 <= data_in;
	if (addr_selector[5]&addr_selector[15])
		data_out <= r_5_15;
		if (write_en==1'b1)
			r_5_15 <= data_in;
	if (addr_selector[5]&addr_selector[16])
		data_out <= r_5_16;
		if (write_en==1'b1)
			r_5_16 <= data_in;
	if (addr_selector[5]&addr_selector[17])
		data_out <= r_5_17;
		if (write_en==1'b1)
			r_5_17 <= data_in;
	if (addr_selector[5]&addr_selector[18])
		data_out <= r_5_18;
		if (write_en==1'b1)
			r_5_18 <= data_in;
	if (addr_selector[5]&addr_selector[19])
		data_out <= r_5_19;
		if (write_en==1'b1)
			r_5_19 <= data_in;
	if (addr_selector[5]&addr_selector[20])
		data_out <= r_5_20;
		if (write_en==1'b1)
			r_5_20 <= data_in;
	if (addr_selector[5]&addr_selector[21])
		data_out <= r_5_21;
		if (write_en==1'b1)
			r_5_21 <= data_in;
	if (addr_selector[5]&addr_selector[22])
		data_out <= r_5_22;
		if (write_en==1'b1)
			r_5_22 <= data_in;
	if (addr_selector[5]&addr_selector[23])
		data_out <= r_5_23;
		if (write_en==1'b1)
			r_5_23 <= data_in;
	if (addr_selector[5]&addr_selector[24])
		data_out <= r_5_24;
		if (write_en==1'b1)
			r_5_24 <= data_in;
	if (addr_selector[5]&addr_selector[25])
		data_out <= r_5_25;
		if (write_en==1'b1)
			r_5_25 <= data_in;
	if (addr_selector[5]&addr_selector[26])
		data_out <= r_5_26;
		if (write_en==1'b1)
			r_5_26 <= data_in;
	if (addr_selector[5]&addr_selector[27])
		data_out <= r_5_27;
		if (write_en==1'b1)
			r_5_27 <= data_in;
	if (addr_selector[5]&addr_selector[28])
		data_out <= r_5_28;
		if (write_en==1'b1)
			r_5_28 <= data_in;
	if (addr_selector[5]&addr_selector[29])
		data_out <= r_5_29;
		if (write_en==1'b1)
			r_5_29 <= data_in;
	if (addr_selector[5]&addr_selector[30])
		data_out <= r_5_30;
		if (write_en==1'b1)
			r_5_30 <= data_in;
	if (addr_selector[5]&addr_selector[31])
		data_out <= r_5_31;
		if (write_en==1'b1)
			r_5_31 <= data_in;
	if (addr_selector[5]&addr_selector[32])
		data_out <= r_5_32;
		if (write_en==1'b1)
			r_5_32 <= data_in;
	if (addr_selector[5]&addr_selector[33])
		data_out <= r_5_33;
		if (write_en==1'b1)
			r_5_33 <= data_in;
	if (addr_selector[5]&addr_selector[34])
		data_out <= r_5_34;
		if (write_en==1'b1)
			r_5_34 <= data_in;
	if (addr_selector[5]&addr_selector[35])
		data_out <= r_5_35;
		if (write_en==1'b1)
			r_5_35 <= data_in;
	if (addr_selector[5]&addr_selector[36])
		data_out <= r_5_36;
		if (write_en==1'b1)
			r_5_36 <= data_in;
	if (addr_selector[5]&addr_selector[37])
		data_out <= r_5_37;
		if (write_en==1'b1)
			r_5_37 <= data_in;
	if (addr_selector[5]&addr_selector[38])
		data_out <= r_5_38;
		if (write_en==1'b1)
			r_5_38 <= data_in;
	if (addr_selector[5]&addr_selector[39])
		data_out <= r_5_39;
		if (write_en==1'b1)
			r_5_39 <= data_in;
	if (addr_selector[5]&addr_selector[40])
		data_out <= r_5_40;
		if (write_en==1'b1)
			r_5_40 <= data_in;
	if (addr_selector[5]&addr_selector[41])
		data_out <= r_5_41;
		if (write_en==1'b1)
			r_5_41 <= data_in;
	if (addr_selector[5]&addr_selector[42])
		data_out <= r_5_42;
		if (write_en==1'b1)
			r_5_42 <= data_in;
	if (addr_selector[5]&addr_selector[43])
		data_out <= r_5_43;
		if (write_en==1'b1)
			r_5_43 <= data_in;
	if (addr_selector[5]&addr_selector[44])
		data_out <= r_5_44;
		if (write_en==1'b1)
			r_5_44 <= data_in;
	if (addr_selector[5]&addr_selector[45])
		data_out <= r_5_45;
		if (write_en==1'b1)
			r_5_45 <= data_in;
	if (addr_selector[5]&addr_selector[46])
		data_out <= r_5_46;
		if (write_en==1'b1)
			r_5_46 <= data_in;
	if (addr_selector[5]&addr_selector[47])
		data_out <= r_5_47;
		if (write_en==1'b1)
			r_5_47 <= data_in;
	if (addr_selector[5]&addr_selector[48])
		data_out <= r_5_48;
		if (write_en==1'b1)
			r_5_48 <= data_in;
	if (addr_selector[5]&addr_selector[49])
		data_out <= r_5_49;
		if (write_en==1'b1)
			r_5_49 <= data_in;
	if (addr_selector[5]&addr_selector[50])
		data_out <= r_5_50;
		if (write_en==1'b1)
			r_5_50 <= data_in;
	if (addr_selector[5]&addr_selector[51])
		data_out <= r_5_51;
		if (write_en==1'b1)
			r_5_51 <= data_in;
	if (addr_selector[5]&addr_selector[52])
		data_out <= r_5_52;
		if (write_en==1'b1)
			r_5_52 <= data_in;
	if (addr_selector[5]&addr_selector[53])
		data_out <= r_5_53;
		if (write_en==1'b1)
			r_5_53 <= data_in;
	if (addr_selector[5]&addr_selector[54])
		data_out <= r_5_54;
		if (write_en==1'b1)
			r_5_54 <= data_in;
	if (addr_selector[5]&addr_selector[55])
		data_out <= r_5_55;
		if (write_en==1'b1)
			r_5_55 <= data_in;
	if (addr_selector[5]&addr_selector[56])
		data_out <= r_5_56;
		if (write_en==1'b1)
			r_5_56 <= data_in;
	if (addr_selector[5]&addr_selector[57])
		data_out <= r_5_57;
		if (write_en==1'b1)
			r_5_57 <= data_in;
	if (addr_selector[5]&addr_selector[58])
		data_out <= r_5_58;
		if (write_en==1'b1)
			r_5_58 <= data_in;
	if (addr_selector[5]&addr_selector[59])
		data_out <= r_5_59;
		if (write_en==1'b1)
			r_5_59 <= data_in;
	if (addr_selector[5]&addr_selector[60])
		data_out <= r_5_60;
		if (write_en==1'b1)
			r_5_60 <= data_in;
	if (addr_selector[5]&addr_selector[61])
		data_out <= r_5_61;
		if (write_en==1'b1)
			r_5_61 <= data_in;
	if (addr_selector[5]&addr_selector[62])
		data_out <= r_5_62;
		if (write_en==1'b1)
			r_5_62 <= data_in;
	if (addr_selector[5]&addr_selector[63])
		data_out <= r_5_63;
		if (write_en==1'b1)
			r_5_63 <= data_in;
	if (addr_selector[6]&addr_selector[0])
		data_out <= r_6_0;
		if (write_en==1'b1)
			r_6_0 <= data_in;
	if (addr_selector[6]&addr_selector[1])
		data_out <= r_6_1;
		if (write_en==1'b1)
			r_6_1 <= data_in;
	if (addr_selector[6]&addr_selector[2])
		data_out <= r_6_2;
		if (write_en==1'b1)
			r_6_2 <= data_in;
	if (addr_selector[6]&addr_selector[3])
		data_out <= r_6_3;
		if (write_en==1'b1)
			r_6_3 <= data_in;
	if (addr_selector[6]&addr_selector[4])
		data_out <= r_6_4;
		if (write_en==1'b1)
			r_6_4 <= data_in;
	if (addr_selector[6]&addr_selector[5])
		data_out <= r_6_5;
		if (write_en==1'b1)
			r_6_5 <= data_in;
	if (addr_selector[6]&addr_selector[6])
		data_out <= r_6_6;
		if (write_en==1'b1)
			r_6_6 <= data_in;
	if (addr_selector[6]&addr_selector[7])
		data_out <= r_6_7;
		if (write_en==1'b1)
			r_6_7 <= data_in;
	if (addr_selector[6]&addr_selector[8])
		data_out <= r_6_8;
		if (write_en==1'b1)
			r_6_8 <= data_in;
	if (addr_selector[6]&addr_selector[9])
		data_out <= r_6_9;
		if (write_en==1'b1)
			r_6_9 <= data_in;
	if (addr_selector[6]&addr_selector[10])
		data_out <= r_6_10;
		if (write_en==1'b1)
			r_6_10 <= data_in;
	if (addr_selector[6]&addr_selector[11])
		data_out <= r_6_11;
		if (write_en==1'b1)
			r_6_11 <= data_in;
	if (addr_selector[6]&addr_selector[12])
		data_out <= r_6_12;
		if (write_en==1'b1)
			r_6_12 <= data_in;
	if (addr_selector[6]&addr_selector[13])
		data_out <= r_6_13;
		if (write_en==1'b1)
			r_6_13 <= data_in;
	if (addr_selector[6]&addr_selector[14])
		data_out <= r_6_14;
		if (write_en==1'b1)
			r_6_14 <= data_in;
	if (addr_selector[6]&addr_selector[15])
		data_out <= r_6_15;
		if (write_en==1'b1)
			r_6_15 <= data_in;
	if (addr_selector[6]&addr_selector[16])
		data_out <= r_6_16;
		if (write_en==1'b1)
			r_6_16 <= data_in;
	if (addr_selector[6]&addr_selector[17])
		data_out <= r_6_17;
		if (write_en==1'b1)
			r_6_17 <= data_in;
	if (addr_selector[6]&addr_selector[18])
		data_out <= r_6_18;
		if (write_en==1'b1)
			r_6_18 <= data_in;
	if (addr_selector[6]&addr_selector[19])
		data_out <= r_6_19;
		if (write_en==1'b1)
			r_6_19 <= data_in;
	if (addr_selector[6]&addr_selector[20])
		data_out <= r_6_20;
		if (write_en==1'b1)
			r_6_20 <= data_in;
	if (addr_selector[6]&addr_selector[21])
		data_out <= r_6_21;
		if (write_en==1'b1)
			r_6_21 <= data_in;
	if (addr_selector[6]&addr_selector[22])
		data_out <= r_6_22;
		if (write_en==1'b1)
			r_6_22 <= data_in;
	if (addr_selector[6]&addr_selector[23])
		data_out <= r_6_23;
		if (write_en==1'b1)
			r_6_23 <= data_in;
	if (addr_selector[6]&addr_selector[24])
		data_out <= r_6_24;
		if (write_en==1'b1)
			r_6_24 <= data_in;
	if (addr_selector[6]&addr_selector[25])
		data_out <= r_6_25;
		if (write_en==1'b1)
			r_6_25 <= data_in;
	if (addr_selector[6]&addr_selector[26])
		data_out <= r_6_26;
		if (write_en==1'b1)
			r_6_26 <= data_in;
	if (addr_selector[6]&addr_selector[27])
		data_out <= r_6_27;
		if (write_en==1'b1)
			r_6_27 <= data_in;
	if (addr_selector[6]&addr_selector[28])
		data_out <= r_6_28;
		if (write_en==1'b1)
			r_6_28 <= data_in;
	if (addr_selector[6]&addr_selector[29])
		data_out <= r_6_29;
		if (write_en==1'b1)
			r_6_29 <= data_in;
	if (addr_selector[6]&addr_selector[30])
		data_out <= r_6_30;
		if (write_en==1'b1)
			r_6_30 <= data_in;
	if (addr_selector[6]&addr_selector[31])
		data_out <= r_6_31;
		if (write_en==1'b1)
			r_6_31 <= data_in;
	if (addr_selector[6]&addr_selector[32])
		data_out <= r_6_32;
		if (write_en==1'b1)
			r_6_32 <= data_in;
	if (addr_selector[6]&addr_selector[33])
		data_out <= r_6_33;
		if (write_en==1'b1)
			r_6_33 <= data_in;
	if (addr_selector[6]&addr_selector[34])
		data_out <= r_6_34;
		if (write_en==1'b1)
			r_6_34 <= data_in;
	if (addr_selector[6]&addr_selector[35])
		data_out <= r_6_35;
		if (write_en==1'b1)
			r_6_35 <= data_in;
	if (addr_selector[6]&addr_selector[36])
		data_out <= r_6_36;
		if (write_en==1'b1)
			r_6_36 <= data_in;
	if (addr_selector[6]&addr_selector[37])
		data_out <= r_6_37;
		if (write_en==1'b1)
			r_6_37 <= data_in;
	if (addr_selector[6]&addr_selector[38])
		data_out <= r_6_38;
		if (write_en==1'b1)
			r_6_38 <= data_in;
	if (addr_selector[6]&addr_selector[39])
		data_out <= r_6_39;
		if (write_en==1'b1)
			r_6_39 <= data_in;
	if (addr_selector[6]&addr_selector[40])
		data_out <= r_6_40;
		if (write_en==1'b1)
			r_6_40 <= data_in;
	if (addr_selector[6]&addr_selector[41])
		data_out <= r_6_41;
		if (write_en==1'b1)
			r_6_41 <= data_in;
	if (addr_selector[6]&addr_selector[42])
		data_out <= r_6_42;
		if (write_en==1'b1)
			r_6_42 <= data_in;
	if (addr_selector[6]&addr_selector[43])
		data_out <= r_6_43;
		if (write_en==1'b1)
			r_6_43 <= data_in;
	if (addr_selector[6]&addr_selector[44])
		data_out <= r_6_44;
		if (write_en==1'b1)
			r_6_44 <= data_in;
	if (addr_selector[6]&addr_selector[45])
		data_out <= r_6_45;
		if (write_en==1'b1)
			r_6_45 <= data_in;
	if (addr_selector[6]&addr_selector[46])
		data_out <= r_6_46;
		if (write_en==1'b1)
			r_6_46 <= data_in;
	if (addr_selector[6]&addr_selector[47])
		data_out <= r_6_47;
		if (write_en==1'b1)
			r_6_47 <= data_in;
	if (addr_selector[6]&addr_selector[48])
		data_out <= r_6_48;
		if (write_en==1'b1)
			r_6_48 <= data_in;
	if (addr_selector[6]&addr_selector[49])
		data_out <= r_6_49;
		if (write_en==1'b1)
			r_6_49 <= data_in;
	if (addr_selector[6]&addr_selector[50])
		data_out <= r_6_50;
		if (write_en==1'b1)
			r_6_50 <= data_in;
	if (addr_selector[6]&addr_selector[51])
		data_out <= r_6_51;
		if (write_en==1'b1)
			r_6_51 <= data_in;
	if (addr_selector[6]&addr_selector[52])
		data_out <= r_6_52;
		if (write_en==1'b1)
			r_6_52 <= data_in;
	if (addr_selector[6]&addr_selector[53])
		data_out <= r_6_53;
		if (write_en==1'b1)
			r_6_53 <= data_in;
	if (addr_selector[6]&addr_selector[54])
		data_out <= r_6_54;
		if (write_en==1'b1)
			r_6_54 <= data_in;
	if (addr_selector[6]&addr_selector[55])
		data_out <= r_6_55;
		if (write_en==1'b1)
			r_6_55 <= data_in;
	if (addr_selector[6]&addr_selector[56])
		data_out <= r_6_56;
		if (write_en==1'b1)
			r_6_56 <= data_in;
	if (addr_selector[6]&addr_selector[57])
		data_out <= r_6_57;
		if (write_en==1'b1)
			r_6_57 <= data_in;
	if (addr_selector[6]&addr_selector[58])
		data_out <= r_6_58;
		if (write_en==1'b1)
			r_6_58 <= data_in;
	if (addr_selector[6]&addr_selector[59])
		data_out <= r_6_59;
		if (write_en==1'b1)
			r_6_59 <= data_in;
	if (addr_selector[6]&addr_selector[60])
		data_out <= r_6_60;
		if (write_en==1'b1)
			r_6_60 <= data_in;
	if (addr_selector[6]&addr_selector[61])
		data_out <= r_6_61;
		if (write_en==1'b1)
			r_6_61 <= data_in;
	if (addr_selector[6]&addr_selector[62])
		data_out <= r_6_62;
		if (write_en==1'b1)
			r_6_62 <= data_in;
	if (addr_selector[6]&addr_selector[63])
		data_out <= r_6_63;
		if (write_en==1'b1)
			r_6_63 <= data_in;
	if (addr_selector[7]&addr_selector[0])
		data_out <= r_7_0;
		if (write_en==1'b1)
			r_7_0 <= data_in;
	if (addr_selector[7]&addr_selector[1])
		data_out <= r_7_1;
		if (write_en==1'b1)
			r_7_1 <= data_in;
	if (addr_selector[7]&addr_selector[2])
		data_out <= r_7_2;
		if (write_en==1'b1)
			r_7_2 <= data_in;
	if (addr_selector[7]&addr_selector[3])
		data_out <= r_7_3;
		if (write_en==1'b1)
			r_7_3 <= data_in;
	if (addr_selector[7]&addr_selector[4])
		data_out <= r_7_4;
		if (write_en==1'b1)
			r_7_4 <= data_in;
	if (addr_selector[7]&addr_selector[5])
		data_out <= r_7_5;
		if (write_en==1'b1)
			r_7_5 <= data_in;
	if (addr_selector[7]&addr_selector[6])
		data_out <= r_7_6;
		if (write_en==1'b1)
			r_7_6 <= data_in;
	if (addr_selector[7]&addr_selector[7])
		data_out <= r_7_7;
		if (write_en==1'b1)
			r_7_7 <= data_in;
	if (addr_selector[7]&addr_selector[8])
		data_out <= r_7_8;
		if (write_en==1'b1)
			r_7_8 <= data_in;
	if (addr_selector[7]&addr_selector[9])
		data_out <= r_7_9;
		if (write_en==1'b1)
			r_7_9 <= data_in;
	if (addr_selector[7]&addr_selector[10])
		data_out <= r_7_10;
		if (write_en==1'b1)
			r_7_10 <= data_in;
	if (addr_selector[7]&addr_selector[11])
		data_out <= r_7_11;
		if (write_en==1'b1)
			r_7_11 <= data_in;
	if (addr_selector[7]&addr_selector[12])
		data_out <= r_7_12;
		if (write_en==1'b1)
			r_7_12 <= data_in;
	if (addr_selector[7]&addr_selector[13])
		data_out <= r_7_13;
		if (write_en==1'b1)
			r_7_13 <= data_in;
	if (addr_selector[7]&addr_selector[14])
		data_out <= r_7_14;
		if (write_en==1'b1)
			r_7_14 <= data_in;
	if (addr_selector[7]&addr_selector[15])
		data_out <= r_7_15;
		if (write_en==1'b1)
			r_7_15 <= data_in;
	if (addr_selector[7]&addr_selector[16])
		data_out <= r_7_16;
		if (write_en==1'b1)
			r_7_16 <= data_in;
	if (addr_selector[7]&addr_selector[17])
		data_out <= r_7_17;
		if (write_en==1'b1)
			r_7_17 <= data_in;
	if (addr_selector[7]&addr_selector[18])
		data_out <= r_7_18;
		if (write_en==1'b1)
			r_7_18 <= data_in;
	if (addr_selector[7]&addr_selector[19])
		data_out <= r_7_19;
		if (write_en==1'b1)
			r_7_19 <= data_in;
	if (addr_selector[7]&addr_selector[20])
		data_out <= r_7_20;
		if (write_en==1'b1)
			r_7_20 <= data_in;
	if (addr_selector[7]&addr_selector[21])
		data_out <= r_7_21;
		if (write_en==1'b1)
			r_7_21 <= data_in;
	if (addr_selector[7]&addr_selector[22])
		data_out <= r_7_22;
		if (write_en==1'b1)
			r_7_22 <= data_in;
	if (addr_selector[7]&addr_selector[23])
		data_out <= r_7_23;
		if (write_en==1'b1)
			r_7_23 <= data_in;
	if (addr_selector[7]&addr_selector[24])
		data_out <= r_7_24;
		if (write_en==1'b1)
			r_7_24 <= data_in;
	if (addr_selector[7]&addr_selector[25])
		data_out <= r_7_25;
		if (write_en==1'b1)
			r_7_25 <= data_in;
	if (addr_selector[7]&addr_selector[26])
		data_out <= r_7_26;
		if (write_en==1'b1)
			r_7_26 <= data_in;
	if (addr_selector[7]&addr_selector[27])
		data_out <= r_7_27;
		if (write_en==1'b1)
			r_7_27 <= data_in;
	if (addr_selector[7]&addr_selector[28])
		data_out <= r_7_28;
		if (write_en==1'b1)
			r_7_28 <= data_in;
	if (addr_selector[7]&addr_selector[29])
		data_out <= r_7_29;
		if (write_en==1'b1)
			r_7_29 <= data_in;
	if (addr_selector[7]&addr_selector[30])
		data_out <= r_7_30;
		if (write_en==1'b1)
			r_7_30 <= data_in;
	if (addr_selector[7]&addr_selector[31])
		data_out <= r_7_31;
		if (write_en==1'b1)
			r_7_31 <= data_in;
	if (addr_selector[7]&addr_selector[32])
		data_out <= r_7_32;
		if (write_en==1'b1)
			r_7_32 <= data_in;
	if (addr_selector[7]&addr_selector[33])
		data_out <= r_7_33;
		if (write_en==1'b1)
			r_7_33 <= data_in;
	if (addr_selector[7]&addr_selector[34])
		data_out <= r_7_34;
		if (write_en==1'b1)
			r_7_34 <= data_in;
	if (addr_selector[7]&addr_selector[35])
		data_out <= r_7_35;
		if (write_en==1'b1)
			r_7_35 <= data_in;
	if (addr_selector[7]&addr_selector[36])
		data_out <= r_7_36;
		if (write_en==1'b1)
			r_7_36 <= data_in;
	if (addr_selector[7]&addr_selector[37])
		data_out <= r_7_37;
		if (write_en==1'b1)
			r_7_37 <= data_in;
	if (addr_selector[7]&addr_selector[38])
		data_out <= r_7_38;
		if (write_en==1'b1)
			r_7_38 <= data_in;
	if (addr_selector[7]&addr_selector[39])
		data_out <= r_7_39;
		if (write_en==1'b1)
			r_7_39 <= data_in;
	if (addr_selector[7]&addr_selector[40])
		data_out <= r_7_40;
		if (write_en==1'b1)
			r_7_40 <= data_in;
	if (addr_selector[7]&addr_selector[41])
		data_out <= r_7_41;
		if (write_en==1'b1)
			r_7_41 <= data_in;
	if (addr_selector[7]&addr_selector[42])
		data_out <= r_7_42;
		if (write_en==1'b1)
			r_7_42 <= data_in;
	if (addr_selector[7]&addr_selector[43])
		data_out <= r_7_43;
		if (write_en==1'b1)
			r_7_43 <= data_in;
	if (addr_selector[7]&addr_selector[44])
		data_out <= r_7_44;
		if (write_en==1'b1)
			r_7_44 <= data_in;
	if (addr_selector[7]&addr_selector[45])
		data_out <= r_7_45;
		if (write_en==1'b1)
			r_7_45 <= data_in;
	if (addr_selector[7]&addr_selector[46])
		data_out <= r_7_46;
		if (write_en==1'b1)
			r_7_46 <= data_in;
	if (addr_selector[7]&addr_selector[47])
		data_out <= r_7_47;
		if (write_en==1'b1)
			r_7_47 <= data_in;
	if (addr_selector[7]&addr_selector[48])
		data_out <= r_7_48;
		if (write_en==1'b1)
			r_7_48 <= data_in;
	if (addr_selector[7]&addr_selector[49])
		data_out <= r_7_49;
		if (write_en==1'b1)
			r_7_49 <= data_in;
	if (addr_selector[7]&addr_selector[50])
		data_out <= r_7_50;
		if (write_en==1'b1)
			r_7_50 <= data_in;
	if (addr_selector[7]&addr_selector[51])
		data_out <= r_7_51;
		if (write_en==1'b1)
			r_7_51 <= data_in;
	if (addr_selector[7]&addr_selector[52])
		data_out <= r_7_52;
		if (write_en==1'b1)
			r_7_52 <= data_in;
	if (addr_selector[7]&addr_selector[53])
		data_out <= r_7_53;
		if (write_en==1'b1)
			r_7_53 <= data_in;
	if (addr_selector[7]&addr_selector[54])
		data_out <= r_7_54;
		if (write_en==1'b1)
			r_7_54 <= data_in;
	if (addr_selector[7]&addr_selector[55])
		data_out <= r_7_55;
		if (write_en==1'b1)
			r_7_55 <= data_in;
	if (addr_selector[7]&addr_selector[56])
		data_out <= r_7_56;
		if (write_en==1'b1)
			r_7_56 <= data_in;
	if (addr_selector[7]&addr_selector[57])
		data_out <= r_7_57;
		if (write_en==1'b1)
			r_7_57 <= data_in;
	if (addr_selector[7]&addr_selector[58])
		data_out <= r_7_58;
		if (write_en==1'b1)
			r_7_58 <= data_in;
	if (addr_selector[7]&addr_selector[59])
		data_out <= r_7_59;
		if (write_en==1'b1)
			r_7_59 <= data_in;
	if (addr_selector[7]&addr_selector[60])
		data_out <= r_7_60;
		if (write_en==1'b1)
			r_7_60 <= data_in;
	if (addr_selector[7]&addr_selector[61])
		data_out <= r_7_61;
		if (write_en==1'b1)
			r_7_61 <= data_in;
	if (addr_selector[7]&addr_selector[62])
		data_out <= r_7_62;
		if (write_en==1'b1)
			r_7_62 <= data_in;
	if (addr_selector[7]&addr_selector[63])
		data_out <= r_7_63;
		if (write_en==1'b1)
			r_7_63 <= data_in;
	if (addr_selector[8]&addr_selector[0])
		data_out <= r_8_0;
		if (write_en==1'b1)
			r_8_0 <= data_in;
	if (addr_selector[8]&addr_selector[1])
		data_out <= r_8_1;
		if (write_en==1'b1)
			r_8_1 <= data_in;
	if (addr_selector[8]&addr_selector[2])
		data_out <= r_8_2;
		if (write_en==1'b1)
			r_8_2 <= data_in;
	if (addr_selector[8]&addr_selector[3])
		data_out <= r_8_3;
		if (write_en==1'b1)
			r_8_3 <= data_in;
	if (addr_selector[8]&addr_selector[4])
		data_out <= r_8_4;
		if (write_en==1'b1)
			r_8_4 <= data_in;
	if (addr_selector[8]&addr_selector[5])
		data_out <= r_8_5;
		if (write_en==1'b1)
			r_8_5 <= data_in;
	if (addr_selector[8]&addr_selector[6])
		data_out <= r_8_6;
		if (write_en==1'b1)
			r_8_6 <= data_in;
	if (addr_selector[8]&addr_selector[7])
		data_out <= r_8_7;
		if (write_en==1'b1)
			r_8_7 <= data_in;
	if (addr_selector[8]&addr_selector[8])
		data_out <= r_8_8;
		if (write_en==1'b1)
			r_8_8 <= data_in;
	if (addr_selector[8]&addr_selector[9])
		data_out <= r_8_9;
		if (write_en==1'b1)
			r_8_9 <= data_in;
	if (addr_selector[8]&addr_selector[10])
		data_out <= r_8_10;
		if (write_en==1'b1)
			r_8_10 <= data_in;
	if (addr_selector[8]&addr_selector[11])
		data_out <= r_8_11;
		if (write_en==1'b1)
			r_8_11 <= data_in;
	if (addr_selector[8]&addr_selector[12])
		data_out <= r_8_12;
		if (write_en==1'b1)
			r_8_12 <= data_in;
	if (addr_selector[8]&addr_selector[13])
		data_out <= r_8_13;
		if (write_en==1'b1)
			r_8_13 <= data_in;
	if (addr_selector[8]&addr_selector[14])
		data_out <= r_8_14;
		if (write_en==1'b1)
			r_8_14 <= data_in;
	if (addr_selector[8]&addr_selector[15])
		data_out <= r_8_15;
		if (write_en==1'b1)
			r_8_15 <= data_in;
	if (addr_selector[8]&addr_selector[16])
		data_out <= r_8_16;
		if (write_en==1'b1)
			r_8_16 <= data_in;
	if (addr_selector[8]&addr_selector[17])
		data_out <= r_8_17;
		if (write_en==1'b1)
			r_8_17 <= data_in;
	if (addr_selector[8]&addr_selector[18])
		data_out <= r_8_18;
		if (write_en==1'b1)
			r_8_18 <= data_in;
	if (addr_selector[8]&addr_selector[19])
		data_out <= r_8_19;
		if (write_en==1'b1)
			r_8_19 <= data_in;
	if (addr_selector[8]&addr_selector[20])
		data_out <= r_8_20;
		if (write_en==1'b1)
			r_8_20 <= data_in;
	if (addr_selector[8]&addr_selector[21])
		data_out <= r_8_21;
		if (write_en==1'b1)
			r_8_21 <= data_in;
	if (addr_selector[8]&addr_selector[22])
		data_out <= r_8_22;
		if (write_en==1'b1)
			r_8_22 <= data_in;
	if (addr_selector[8]&addr_selector[23])
		data_out <= r_8_23;
		if (write_en==1'b1)
			r_8_23 <= data_in;
	if (addr_selector[8]&addr_selector[24])
		data_out <= r_8_24;
		if (write_en==1'b1)
			r_8_24 <= data_in;
	if (addr_selector[8]&addr_selector[25])
		data_out <= r_8_25;
		if (write_en==1'b1)
			r_8_25 <= data_in;
	if (addr_selector[8]&addr_selector[26])
		data_out <= r_8_26;
		if (write_en==1'b1)
			r_8_26 <= data_in;
	if (addr_selector[8]&addr_selector[27])
		data_out <= r_8_27;
		if (write_en==1'b1)
			r_8_27 <= data_in;
	if (addr_selector[8]&addr_selector[28])
		data_out <= r_8_28;
		if (write_en==1'b1)
			r_8_28 <= data_in;
	if (addr_selector[8]&addr_selector[29])
		data_out <= r_8_29;
		if (write_en==1'b1)
			r_8_29 <= data_in;
	if (addr_selector[8]&addr_selector[30])
		data_out <= r_8_30;
		if (write_en==1'b1)
			r_8_30 <= data_in;
	if (addr_selector[8]&addr_selector[31])
		data_out <= r_8_31;
		if (write_en==1'b1)
			r_8_31 <= data_in;
	if (addr_selector[8]&addr_selector[32])
		data_out <= r_8_32;
		if (write_en==1'b1)
			r_8_32 <= data_in;
	if (addr_selector[8]&addr_selector[33])
		data_out <= r_8_33;
		if (write_en==1'b1)
			r_8_33 <= data_in;
	if (addr_selector[8]&addr_selector[34])
		data_out <= r_8_34;
		if (write_en==1'b1)
			r_8_34 <= data_in;
	if (addr_selector[8]&addr_selector[35])
		data_out <= r_8_35;
		if (write_en==1'b1)
			r_8_35 <= data_in;
	if (addr_selector[8]&addr_selector[36])
		data_out <= r_8_36;
		if (write_en==1'b1)
			r_8_36 <= data_in;
	if (addr_selector[8]&addr_selector[37])
		data_out <= r_8_37;
		if (write_en==1'b1)
			r_8_37 <= data_in;
	if (addr_selector[8]&addr_selector[38])
		data_out <= r_8_38;
		if (write_en==1'b1)
			r_8_38 <= data_in;
	if (addr_selector[8]&addr_selector[39])
		data_out <= r_8_39;
		if (write_en==1'b1)
			r_8_39 <= data_in;
	if (addr_selector[8]&addr_selector[40])
		data_out <= r_8_40;
		if (write_en==1'b1)
			r_8_40 <= data_in;
	if (addr_selector[8]&addr_selector[41])
		data_out <= r_8_41;
		if (write_en==1'b1)
			r_8_41 <= data_in;
	if (addr_selector[8]&addr_selector[42])
		data_out <= r_8_42;
		if (write_en==1'b1)
			r_8_42 <= data_in;
	if (addr_selector[8]&addr_selector[43])
		data_out <= r_8_43;
		if (write_en==1'b1)
			r_8_43 <= data_in;
	if (addr_selector[8]&addr_selector[44])
		data_out <= r_8_44;
		if (write_en==1'b1)
			r_8_44 <= data_in;
	if (addr_selector[8]&addr_selector[45])
		data_out <= r_8_45;
		if (write_en==1'b1)
			r_8_45 <= data_in;
	if (addr_selector[8]&addr_selector[46])
		data_out <= r_8_46;
		if (write_en==1'b1)
			r_8_46 <= data_in;
	if (addr_selector[8]&addr_selector[47])
		data_out <= r_8_47;
		if (write_en==1'b1)
			r_8_47 <= data_in;
	if (addr_selector[8]&addr_selector[48])
		data_out <= r_8_48;
		if (write_en==1'b1)
			r_8_48 <= data_in;
	if (addr_selector[8]&addr_selector[49])
		data_out <= r_8_49;
		if (write_en==1'b1)
			r_8_49 <= data_in;
	if (addr_selector[8]&addr_selector[50])
		data_out <= r_8_50;
		if (write_en==1'b1)
			r_8_50 <= data_in;
	if (addr_selector[8]&addr_selector[51])
		data_out <= r_8_51;
		if (write_en==1'b1)
			r_8_51 <= data_in;
	if (addr_selector[8]&addr_selector[52])
		data_out <= r_8_52;
		if (write_en==1'b1)
			r_8_52 <= data_in;
	if (addr_selector[8]&addr_selector[53])
		data_out <= r_8_53;
		if (write_en==1'b1)
			r_8_53 <= data_in;
	if (addr_selector[8]&addr_selector[54])
		data_out <= r_8_54;
		if (write_en==1'b1)
			r_8_54 <= data_in;
	if (addr_selector[8]&addr_selector[55])
		data_out <= r_8_55;
		if (write_en==1'b1)
			r_8_55 <= data_in;
	if (addr_selector[8]&addr_selector[56])
		data_out <= r_8_56;
		if (write_en==1'b1)
			r_8_56 <= data_in;
	if (addr_selector[8]&addr_selector[57])
		data_out <= r_8_57;
		if (write_en==1'b1)
			r_8_57 <= data_in;
	if (addr_selector[8]&addr_selector[58])
		data_out <= r_8_58;
		if (write_en==1'b1)
			r_8_58 <= data_in;
	if (addr_selector[8]&addr_selector[59])
		data_out <= r_8_59;
		if (write_en==1'b1)
			r_8_59 <= data_in;
	if (addr_selector[8]&addr_selector[60])
		data_out <= r_8_60;
		if (write_en==1'b1)
			r_8_60 <= data_in;
	if (addr_selector[8]&addr_selector[61])
		data_out <= r_8_61;
		if (write_en==1'b1)
			r_8_61 <= data_in;
	if (addr_selector[8]&addr_selector[62])
		data_out <= r_8_62;
		if (write_en==1'b1)
			r_8_62 <= data_in;
	if (addr_selector[8]&addr_selector[63])
		data_out <= r_8_63;
		if (write_en==1'b1)
			r_8_63 <= data_in;
	if (addr_selector[9]&addr_selector[0])
		data_out <= r_9_0;
		if (write_en==1'b1)
			r_9_0 <= data_in;
	if (addr_selector[9]&addr_selector[1])
		data_out <= r_9_1;
		if (write_en==1'b1)
			r_9_1 <= data_in;
	if (addr_selector[9]&addr_selector[2])
		data_out <= r_9_2;
		if (write_en==1'b1)
			r_9_2 <= data_in;
	if (addr_selector[9]&addr_selector[3])
		data_out <= r_9_3;
		if (write_en==1'b1)
			r_9_3 <= data_in;
	if (addr_selector[9]&addr_selector[4])
		data_out <= r_9_4;
		if (write_en==1'b1)
			r_9_4 <= data_in;
	if (addr_selector[9]&addr_selector[5])
		data_out <= r_9_5;
		if (write_en==1'b1)
			r_9_5 <= data_in;
	if (addr_selector[9]&addr_selector[6])
		data_out <= r_9_6;
		if (write_en==1'b1)
			r_9_6 <= data_in;
	if (addr_selector[9]&addr_selector[7])
		data_out <= r_9_7;
		if (write_en==1'b1)
			r_9_7 <= data_in;
	if (addr_selector[9]&addr_selector[8])
		data_out <= r_9_8;
		if (write_en==1'b1)
			r_9_8 <= data_in;
	if (addr_selector[9]&addr_selector[9])
		data_out <= r_9_9;
		if (write_en==1'b1)
			r_9_9 <= data_in;
	if (addr_selector[9]&addr_selector[10])
		data_out <= r_9_10;
		if (write_en==1'b1)
			r_9_10 <= data_in;
	if (addr_selector[9]&addr_selector[11])
		data_out <= r_9_11;
		if (write_en==1'b1)
			r_9_11 <= data_in;
	if (addr_selector[9]&addr_selector[12])
		data_out <= r_9_12;
		if (write_en==1'b1)
			r_9_12 <= data_in;
	if (addr_selector[9]&addr_selector[13])
		data_out <= r_9_13;
		if (write_en==1'b1)
			r_9_13 <= data_in;
	if (addr_selector[9]&addr_selector[14])
		data_out <= r_9_14;
		if (write_en==1'b1)
			r_9_14 <= data_in;
	if (addr_selector[9]&addr_selector[15])
		data_out <= r_9_15;
		if (write_en==1'b1)
			r_9_15 <= data_in;
	if (addr_selector[9]&addr_selector[16])
		data_out <= r_9_16;
		if (write_en==1'b1)
			r_9_16 <= data_in;
	if (addr_selector[9]&addr_selector[17])
		data_out <= r_9_17;
		if (write_en==1'b1)
			r_9_17 <= data_in;
	if (addr_selector[9]&addr_selector[18])
		data_out <= r_9_18;
		if (write_en==1'b1)
			r_9_18 <= data_in;
	if (addr_selector[9]&addr_selector[19])
		data_out <= r_9_19;
		if (write_en==1'b1)
			r_9_19 <= data_in;
	if (addr_selector[9]&addr_selector[20])
		data_out <= r_9_20;
		if (write_en==1'b1)
			r_9_20 <= data_in;
	if (addr_selector[9]&addr_selector[21])
		data_out <= r_9_21;
		if (write_en==1'b1)
			r_9_21 <= data_in;
	if (addr_selector[9]&addr_selector[22])
		data_out <= r_9_22;
		if (write_en==1'b1)
			r_9_22 <= data_in;
	if (addr_selector[9]&addr_selector[23])
		data_out <= r_9_23;
		if (write_en==1'b1)
			r_9_23 <= data_in;
	if (addr_selector[9]&addr_selector[24])
		data_out <= r_9_24;
		if (write_en==1'b1)
			r_9_24 <= data_in;
	if (addr_selector[9]&addr_selector[25])
		data_out <= r_9_25;
		if (write_en==1'b1)
			r_9_25 <= data_in;
	if (addr_selector[9]&addr_selector[26])
		data_out <= r_9_26;
		if (write_en==1'b1)
			r_9_26 <= data_in;
	if (addr_selector[9]&addr_selector[27])
		data_out <= r_9_27;
		if (write_en==1'b1)
			r_9_27 <= data_in;
	if (addr_selector[9]&addr_selector[28])
		data_out <= r_9_28;
		if (write_en==1'b1)
			r_9_28 <= data_in;
	if (addr_selector[9]&addr_selector[29])
		data_out <= r_9_29;
		if (write_en==1'b1)
			r_9_29 <= data_in;
	if (addr_selector[9]&addr_selector[30])
		data_out <= r_9_30;
		if (write_en==1'b1)
			r_9_30 <= data_in;
	if (addr_selector[9]&addr_selector[31])
		data_out <= r_9_31;
		if (write_en==1'b1)
			r_9_31 <= data_in;
	if (addr_selector[9]&addr_selector[32])
		data_out <= r_9_32;
		if (write_en==1'b1)
			r_9_32 <= data_in;
	if (addr_selector[9]&addr_selector[33])
		data_out <= r_9_33;
		if (write_en==1'b1)
			r_9_33 <= data_in;
	if (addr_selector[9]&addr_selector[34])
		data_out <= r_9_34;
		if (write_en==1'b1)
			r_9_34 <= data_in;
	if (addr_selector[9]&addr_selector[35])
		data_out <= r_9_35;
		if (write_en==1'b1)
			r_9_35 <= data_in;
	if (addr_selector[9]&addr_selector[36])
		data_out <= r_9_36;
		if (write_en==1'b1)
			r_9_36 <= data_in;
	if (addr_selector[9]&addr_selector[37])
		data_out <= r_9_37;
		if (write_en==1'b1)
			r_9_37 <= data_in;
	if (addr_selector[9]&addr_selector[38])
		data_out <= r_9_38;
		if (write_en==1'b1)
			r_9_38 <= data_in;
	if (addr_selector[9]&addr_selector[39])
		data_out <= r_9_39;
		if (write_en==1'b1)
			r_9_39 <= data_in;
	if (addr_selector[9]&addr_selector[40])
		data_out <= r_9_40;
		if (write_en==1'b1)
			r_9_40 <= data_in;
	if (addr_selector[9]&addr_selector[41])
		data_out <= r_9_41;
		if (write_en==1'b1)
			r_9_41 <= data_in;
	if (addr_selector[9]&addr_selector[42])
		data_out <= r_9_42;
		if (write_en==1'b1)
			r_9_42 <= data_in;
	if (addr_selector[9]&addr_selector[43])
		data_out <= r_9_43;
		if (write_en==1'b1)
			r_9_43 <= data_in;
	if (addr_selector[9]&addr_selector[44])
		data_out <= r_9_44;
		if (write_en==1'b1)
			r_9_44 <= data_in;
	if (addr_selector[9]&addr_selector[45])
		data_out <= r_9_45;
		if (write_en==1'b1)
			r_9_45 <= data_in;
	if (addr_selector[9]&addr_selector[46])
		data_out <= r_9_46;
		if (write_en==1'b1)
			r_9_46 <= data_in;
	if (addr_selector[9]&addr_selector[47])
		data_out <= r_9_47;
		if (write_en==1'b1)
			r_9_47 <= data_in;
	if (addr_selector[9]&addr_selector[48])
		data_out <= r_9_48;
		if (write_en==1'b1)
			r_9_48 <= data_in;
	if (addr_selector[9]&addr_selector[49])
		data_out <= r_9_49;
		if (write_en==1'b1)
			r_9_49 <= data_in;
	if (addr_selector[9]&addr_selector[50])
		data_out <= r_9_50;
		if (write_en==1'b1)
			r_9_50 <= data_in;
	if (addr_selector[9]&addr_selector[51])
		data_out <= r_9_51;
		if (write_en==1'b1)
			r_9_51 <= data_in;
	if (addr_selector[9]&addr_selector[52])
		data_out <= r_9_52;
		if (write_en==1'b1)
			r_9_52 <= data_in;
	if (addr_selector[9]&addr_selector[53])
		data_out <= r_9_53;
		if (write_en==1'b1)
			r_9_53 <= data_in;
	if (addr_selector[9]&addr_selector[54])
		data_out <= r_9_54;
		if (write_en==1'b1)
			r_9_54 <= data_in;
	if (addr_selector[9]&addr_selector[55])
		data_out <= r_9_55;
		if (write_en==1'b1)
			r_9_55 <= data_in;
	if (addr_selector[9]&addr_selector[56])
		data_out <= r_9_56;
		if (write_en==1'b1)
			r_9_56 <= data_in;
	if (addr_selector[9]&addr_selector[57])
		data_out <= r_9_57;
		if (write_en==1'b1)
			r_9_57 <= data_in;
	if (addr_selector[9]&addr_selector[58])
		data_out <= r_9_58;
		if (write_en==1'b1)
			r_9_58 <= data_in;
	if (addr_selector[9]&addr_selector[59])
		data_out <= r_9_59;
		if (write_en==1'b1)
			r_9_59 <= data_in;
	if (addr_selector[9]&addr_selector[60])
		data_out <= r_9_60;
		if (write_en==1'b1)
			r_9_60 <= data_in;
	if (addr_selector[9]&addr_selector[61])
		data_out <= r_9_61;
		if (write_en==1'b1)
			r_9_61 <= data_in;
	if (addr_selector[9]&addr_selector[62])
		data_out <= r_9_62;
		if (write_en==1'b1)
			r_9_62 <= data_in;
	if (addr_selector[9]&addr_selector[63])
		data_out <= r_9_63;
		if (write_en==1'b1)
			r_9_63 <= data_in;
	if (addr_selector[10]&addr_selector[0])
		data_out <= r_10_0;
		if (write_en==1'b1)
			r_10_0 <= data_in;
	if (addr_selector[10]&addr_selector[1])
		data_out <= r_10_1;
		if (write_en==1'b1)
			r_10_1 <= data_in;
	if (addr_selector[10]&addr_selector[2])
		data_out <= r_10_2;
		if (write_en==1'b1)
			r_10_2 <= data_in;
	if (addr_selector[10]&addr_selector[3])
		data_out <= r_10_3;
		if (write_en==1'b1)
			r_10_3 <= data_in;
	if (addr_selector[10]&addr_selector[4])
		data_out <= r_10_4;
		if (write_en==1'b1)
			r_10_4 <= data_in;
	if (addr_selector[10]&addr_selector[5])
		data_out <= r_10_5;
		if (write_en==1'b1)
			r_10_5 <= data_in;
	if (addr_selector[10]&addr_selector[6])
		data_out <= r_10_6;
		if (write_en==1'b1)
			r_10_6 <= data_in;
	if (addr_selector[10]&addr_selector[7])
		data_out <= r_10_7;
		if (write_en==1'b1)
			r_10_7 <= data_in;
	if (addr_selector[10]&addr_selector[8])
		data_out <= r_10_8;
		if (write_en==1'b1)
			r_10_8 <= data_in;
	if (addr_selector[10]&addr_selector[9])
		data_out <= r_10_9;
		if (write_en==1'b1)
			r_10_9 <= data_in;
	if (addr_selector[10]&addr_selector[10])
		data_out <= r_10_10;
		if (write_en==1'b1)
			r_10_10 <= data_in;
	if (addr_selector[10]&addr_selector[11])
		data_out <= r_10_11;
		if (write_en==1'b1)
			r_10_11 <= data_in;
	if (addr_selector[10]&addr_selector[12])
		data_out <= r_10_12;
		if (write_en==1'b1)
			r_10_12 <= data_in;
	if (addr_selector[10]&addr_selector[13])
		data_out <= r_10_13;
		if (write_en==1'b1)
			r_10_13 <= data_in;
	if (addr_selector[10]&addr_selector[14])
		data_out <= r_10_14;
		if (write_en==1'b1)
			r_10_14 <= data_in;
	if (addr_selector[10]&addr_selector[15])
		data_out <= r_10_15;
		if (write_en==1'b1)
			r_10_15 <= data_in;
	if (addr_selector[10]&addr_selector[16])
		data_out <= r_10_16;
		if (write_en==1'b1)
			r_10_16 <= data_in;
	if (addr_selector[10]&addr_selector[17])
		data_out <= r_10_17;
		if (write_en==1'b1)
			r_10_17 <= data_in;
	if (addr_selector[10]&addr_selector[18])
		data_out <= r_10_18;
		if (write_en==1'b1)
			r_10_18 <= data_in;
	if (addr_selector[10]&addr_selector[19])
		data_out <= r_10_19;
		if (write_en==1'b1)
			r_10_19 <= data_in;
	if (addr_selector[10]&addr_selector[20])
		data_out <= r_10_20;
		if (write_en==1'b1)
			r_10_20 <= data_in;
	if (addr_selector[10]&addr_selector[21])
		data_out <= r_10_21;
		if (write_en==1'b1)
			r_10_21 <= data_in;
	if (addr_selector[10]&addr_selector[22])
		data_out <= r_10_22;
		if (write_en==1'b1)
			r_10_22 <= data_in;
	if (addr_selector[10]&addr_selector[23])
		data_out <= r_10_23;
		if (write_en==1'b1)
			r_10_23 <= data_in;
	if (addr_selector[10]&addr_selector[24])
		data_out <= r_10_24;
		if (write_en==1'b1)
			r_10_24 <= data_in;
	if (addr_selector[10]&addr_selector[25])
		data_out <= r_10_25;
		if (write_en==1'b1)
			r_10_25 <= data_in;
	if (addr_selector[10]&addr_selector[26])
		data_out <= r_10_26;
		if (write_en==1'b1)
			r_10_26 <= data_in;
	if (addr_selector[10]&addr_selector[27])
		data_out <= r_10_27;
		if (write_en==1'b1)
			r_10_27 <= data_in;
	if (addr_selector[10]&addr_selector[28])
		data_out <= r_10_28;
		if (write_en==1'b1)
			r_10_28 <= data_in;
	if (addr_selector[10]&addr_selector[29])
		data_out <= r_10_29;
		if (write_en==1'b1)
			r_10_29 <= data_in;
	if (addr_selector[10]&addr_selector[30])
		data_out <= r_10_30;
		if (write_en==1'b1)
			r_10_30 <= data_in;
	if (addr_selector[10]&addr_selector[31])
		data_out <= r_10_31;
		if (write_en==1'b1)
			r_10_31 <= data_in;
	if (addr_selector[10]&addr_selector[32])
		data_out <= r_10_32;
		if (write_en==1'b1)
			r_10_32 <= data_in;
	if (addr_selector[10]&addr_selector[33])
		data_out <= r_10_33;
		if (write_en==1'b1)
			r_10_33 <= data_in;
	if (addr_selector[10]&addr_selector[34])
		data_out <= r_10_34;
		if (write_en==1'b1)
			r_10_34 <= data_in;
	if (addr_selector[10]&addr_selector[35])
		data_out <= r_10_35;
		if (write_en==1'b1)
			r_10_35 <= data_in;
	if (addr_selector[10]&addr_selector[36])
		data_out <= r_10_36;
		if (write_en==1'b1)
			r_10_36 <= data_in;
	if (addr_selector[10]&addr_selector[37])
		data_out <= r_10_37;
		if (write_en==1'b1)
			r_10_37 <= data_in;
	if (addr_selector[10]&addr_selector[38])
		data_out <= r_10_38;
		if (write_en==1'b1)
			r_10_38 <= data_in;
	if (addr_selector[10]&addr_selector[39])
		data_out <= r_10_39;
		if (write_en==1'b1)
			r_10_39 <= data_in;
	if (addr_selector[10]&addr_selector[40])
		data_out <= r_10_40;
		if (write_en==1'b1)
			r_10_40 <= data_in;
	if (addr_selector[10]&addr_selector[41])
		data_out <= r_10_41;
		if (write_en==1'b1)
			r_10_41 <= data_in;
	if (addr_selector[10]&addr_selector[42])
		data_out <= r_10_42;
		if (write_en==1'b1)
			r_10_42 <= data_in;
	if (addr_selector[10]&addr_selector[43])
		data_out <= r_10_43;
		if (write_en==1'b1)
			r_10_43 <= data_in;
	if (addr_selector[10]&addr_selector[44])
		data_out <= r_10_44;
		if (write_en==1'b1)
			r_10_44 <= data_in;
	if (addr_selector[10]&addr_selector[45])
		data_out <= r_10_45;
		if (write_en==1'b1)
			r_10_45 <= data_in;
	if (addr_selector[10]&addr_selector[46])
		data_out <= r_10_46;
		if (write_en==1'b1)
			r_10_46 <= data_in;
	if (addr_selector[10]&addr_selector[47])
		data_out <= r_10_47;
		if (write_en==1'b1)
			r_10_47 <= data_in;
	if (addr_selector[10]&addr_selector[48])
		data_out <= r_10_48;
		if (write_en==1'b1)
			r_10_48 <= data_in;
	if (addr_selector[10]&addr_selector[49])
		data_out <= r_10_49;
		if (write_en==1'b1)
			r_10_49 <= data_in;
	if (addr_selector[10]&addr_selector[50])
		data_out <= r_10_50;
		if (write_en==1'b1)
			r_10_50 <= data_in;
	if (addr_selector[10]&addr_selector[51])
		data_out <= r_10_51;
		if (write_en==1'b1)
			r_10_51 <= data_in;
	if (addr_selector[10]&addr_selector[52])
		data_out <= r_10_52;
		if (write_en==1'b1)
			r_10_52 <= data_in;
	if (addr_selector[10]&addr_selector[53])
		data_out <= r_10_53;
		if (write_en==1'b1)
			r_10_53 <= data_in;
	if (addr_selector[10]&addr_selector[54])
		data_out <= r_10_54;
		if (write_en==1'b1)
			r_10_54 <= data_in;
	if (addr_selector[10]&addr_selector[55])
		data_out <= r_10_55;
		if (write_en==1'b1)
			r_10_55 <= data_in;
	if (addr_selector[10]&addr_selector[56])
		data_out <= r_10_56;
		if (write_en==1'b1)
			r_10_56 <= data_in;
	if (addr_selector[10]&addr_selector[57])
		data_out <= r_10_57;
		if (write_en==1'b1)
			r_10_57 <= data_in;
	if (addr_selector[10]&addr_selector[58])
		data_out <= r_10_58;
		if (write_en==1'b1)
			r_10_58 <= data_in;
	if (addr_selector[10]&addr_selector[59])
		data_out <= r_10_59;
		if (write_en==1'b1)
			r_10_59 <= data_in;
	if (addr_selector[10]&addr_selector[60])
		data_out <= r_10_60;
		if (write_en==1'b1)
			r_10_60 <= data_in;
	if (addr_selector[10]&addr_selector[61])
		data_out <= r_10_61;
		if (write_en==1'b1)
			r_10_61 <= data_in;
	if (addr_selector[10]&addr_selector[62])
		data_out <= r_10_62;
		if (write_en==1'b1)
			r_10_62 <= data_in;
	if (addr_selector[10]&addr_selector[63])
		data_out <= r_10_63;
		if (write_en==1'b1)
			r_10_63 <= data_in;
	if (addr_selector[11]&addr_selector[0])
		data_out <= r_11_0;
		if (write_en==1'b1)
			r_11_0 <= data_in;
	if (addr_selector[11]&addr_selector[1])
		data_out <= r_11_1;
		if (write_en==1'b1)
			r_11_1 <= data_in;
	if (addr_selector[11]&addr_selector[2])
		data_out <= r_11_2;
		if (write_en==1'b1)
			r_11_2 <= data_in;
	if (addr_selector[11]&addr_selector[3])
		data_out <= r_11_3;
		if (write_en==1'b1)
			r_11_3 <= data_in;
	if (addr_selector[11]&addr_selector[4])
		data_out <= r_11_4;
		if (write_en==1'b1)
			r_11_4 <= data_in;
	if (addr_selector[11]&addr_selector[5])
		data_out <= r_11_5;
		if (write_en==1'b1)
			r_11_5 <= data_in;
	if (addr_selector[11]&addr_selector[6])
		data_out <= r_11_6;
		if (write_en==1'b1)
			r_11_6 <= data_in;
	if (addr_selector[11]&addr_selector[7])
		data_out <= r_11_7;
		if (write_en==1'b1)
			r_11_7 <= data_in;
	if (addr_selector[11]&addr_selector[8])
		data_out <= r_11_8;
		if (write_en==1'b1)
			r_11_8 <= data_in;
	if (addr_selector[11]&addr_selector[9])
		data_out <= r_11_9;
		if (write_en==1'b1)
			r_11_9 <= data_in;
	if (addr_selector[11]&addr_selector[10])
		data_out <= r_11_10;
		if (write_en==1'b1)
			r_11_10 <= data_in;
	if (addr_selector[11]&addr_selector[11])
		data_out <= r_11_11;
		if (write_en==1'b1)
			r_11_11 <= data_in;
	if (addr_selector[11]&addr_selector[12])
		data_out <= r_11_12;
		if (write_en==1'b1)
			r_11_12 <= data_in;
	if (addr_selector[11]&addr_selector[13])
		data_out <= r_11_13;
		if (write_en==1'b1)
			r_11_13 <= data_in;
	if (addr_selector[11]&addr_selector[14])
		data_out <= r_11_14;
		if (write_en==1'b1)
			r_11_14 <= data_in;
	if (addr_selector[11]&addr_selector[15])
		data_out <= r_11_15;
		if (write_en==1'b1)
			r_11_15 <= data_in;
	if (addr_selector[11]&addr_selector[16])
		data_out <= r_11_16;
		if (write_en==1'b1)
			r_11_16 <= data_in;
	if (addr_selector[11]&addr_selector[17])
		data_out <= r_11_17;
		if (write_en==1'b1)
			r_11_17 <= data_in;
	if (addr_selector[11]&addr_selector[18])
		data_out <= r_11_18;
		if (write_en==1'b1)
			r_11_18 <= data_in;
	if (addr_selector[11]&addr_selector[19])
		data_out <= r_11_19;
		if (write_en==1'b1)
			r_11_19 <= data_in;
	if (addr_selector[11]&addr_selector[20])
		data_out <= r_11_20;
		if (write_en==1'b1)
			r_11_20 <= data_in;
	if (addr_selector[11]&addr_selector[21])
		data_out <= r_11_21;
		if (write_en==1'b1)
			r_11_21 <= data_in;
	if (addr_selector[11]&addr_selector[22])
		data_out <= r_11_22;
		if (write_en==1'b1)
			r_11_22 <= data_in;
	if (addr_selector[11]&addr_selector[23])
		data_out <= r_11_23;
		if (write_en==1'b1)
			r_11_23 <= data_in;
	if (addr_selector[11]&addr_selector[24])
		data_out <= r_11_24;
		if (write_en==1'b1)
			r_11_24 <= data_in;
	if (addr_selector[11]&addr_selector[25])
		data_out <= r_11_25;
		if (write_en==1'b1)
			r_11_25 <= data_in;
	if (addr_selector[11]&addr_selector[26])
		data_out <= r_11_26;
		if (write_en==1'b1)
			r_11_26 <= data_in;
	if (addr_selector[11]&addr_selector[27])
		data_out <= r_11_27;
		if (write_en==1'b1)
			r_11_27 <= data_in;
	if (addr_selector[11]&addr_selector[28])
		data_out <= r_11_28;
		if (write_en==1'b1)
			r_11_28 <= data_in;
	if (addr_selector[11]&addr_selector[29])
		data_out <= r_11_29;
		if (write_en==1'b1)
			r_11_29 <= data_in;
	if (addr_selector[11]&addr_selector[30])
		data_out <= r_11_30;
		if (write_en==1'b1)
			r_11_30 <= data_in;
	if (addr_selector[11]&addr_selector[31])
		data_out <= r_11_31;
		if (write_en==1'b1)
			r_11_31 <= data_in;
	if (addr_selector[11]&addr_selector[32])
		data_out <= r_11_32;
		if (write_en==1'b1)
			r_11_32 <= data_in;
	if (addr_selector[11]&addr_selector[33])
		data_out <= r_11_33;
		if (write_en==1'b1)
			r_11_33 <= data_in;
	if (addr_selector[11]&addr_selector[34])
		data_out <= r_11_34;
		if (write_en==1'b1)
			r_11_34 <= data_in;
	if (addr_selector[11]&addr_selector[35])
		data_out <= r_11_35;
		if (write_en==1'b1)
			r_11_35 <= data_in;
	if (addr_selector[11]&addr_selector[36])
		data_out <= r_11_36;
		if (write_en==1'b1)
			r_11_36 <= data_in;
	if (addr_selector[11]&addr_selector[37])
		data_out <= r_11_37;
		if (write_en==1'b1)
			r_11_37 <= data_in;
	if (addr_selector[11]&addr_selector[38])
		data_out <= r_11_38;
		if (write_en==1'b1)
			r_11_38 <= data_in;
	if (addr_selector[11]&addr_selector[39])
		data_out <= r_11_39;
		if (write_en==1'b1)
			r_11_39 <= data_in;
	if (addr_selector[11]&addr_selector[40])
		data_out <= r_11_40;
		if (write_en==1'b1)
			r_11_40 <= data_in;
	if (addr_selector[11]&addr_selector[41])
		data_out <= r_11_41;
		if (write_en==1'b1)
			r_11_41 <= data_in;
	if (addr_selector[11]&addr_selector[42])
		data_out <= r_11_42;
		if (write_en==1'b1)
			r_11_42 <= data_in;
	if (addr_selector[11]&addr_selector[43])
		data_out <= r_11_43;
		if (write_en==1'b1)
			r_11_43 <= data_in;
	if (addr_selector[11]&addr_selector[44])
		data_out <= r_11_44;
		if (write_en==1'b1)
			r_11_44 <= data_in;
	if (addr_selector[11]&addr_selector[45])
		data_out <= r_11_45;
		if (write_en==1'b1)
			r_11_45 <= data_in;
	if (addr_selector[11]&addr_selector[46])
		data_out <= r_11_46;
		if (write_en==1'b1)
			r_11_46 <= data_in;
	if (addr_selector[11]&addr_selector[47])
		data_out <= r_11_47;
		if (write_en==1'b1)
			r_11_47 <= data_in;
	if (addr_selector[11]&addr_selector[48])
		data_out <= r_11_48;
		if (write_en==1'b1)
			r_11_48 <= data_in;
	if (addr_selector[11]&addr_selector[49])
		data_out <= r_11_49;
		if (write_en==1'b1)
			r_11_49 <= data_in;
	if (addr_selector[11]&addr_selector[50])
		data_out <= r_11_50;
		if (write_en==1'b1)
			r_11_50 <= data_in;
	if (addr_selector[11]&addr_selector[51])
		data_out <= r_11_51;
		if (write_en==1'b1)
			r_11_51 <= data_in;
	if (addr_selector[11]&addr_selector[52])
		data_out <= r_11_52;
		if (write_en==1'b1)
			r_11_52 <= data_in;
	if (addr_selector[11]&addr_selector[53])
		data_out <= r_11_53;
		if (write_en==1'b1)
			r_11_53 <= data_in;
	if (addr_selector[11]&addr_selector[54])
		data_out <= r_11_54;
		if (write_en==1'b1)
			r_11_54 <= data_in;
	if (addr_selector[11]&addr_selector[55])
		data_out <= r_11_55;
		if (write_en==1'b1)
			r_11_55 <= data_in;
	if (addr_selector[11]&addr_selector[56])
		data_out <= r_11_56;
		if (write_en==1'b1)
			r_11_56 <= data_in;
	if (addr_selector[11]&addr_selector[57])
		data_out <= r_11_57;
		if (write_en==1'b1)
			r_11_57 <= data_in;
	if (addr_selector[11]&addr_selector[58])
		data_out <= r_11_58;
		if (write_en==1'b1)
			r_11_58 <= data_in;
	if (addr_selector[11]&addr_selector[59])
		data_out <= r_11_59;
		if (write_en==1'b1)
			r_11_59 <= data_in;
	if (addr_selector[11]&addr_selector[60])
		data_out <= r_11_60;
		if (write_en==1'b1)
			r_11_60 <= data_in;
	if (addr_selector[11]&addr_selector[61])
		data_out <= r_11_61;
		if (write_en==1'b1)
			r_11_61 <= data_in;
	if (addr_selector[11]&addr_selector[62])
		data_out <= r_11_62;
		if (write_en==1'b1)
			r_11_62 <= data_in;
	if (addr_selector[11]&addr_selector[63])
		data_out <= r_11_63;
		if (write_en==1'b1)
			r_11_63 <= data_in;
	if (addr_selector[12]&addr_selector[0])
		data_out <= r_12_0;
		if (write_en==1'b1)
			r_12_0 <= data_in;
	if (addr_selector[12]&addr_selector[1])
		data_out <= r_12_1;
		if (write_en==1'b1)
			r_12_1 <= data_in;
	if (addr_selector[12]&addr_selector[2])
		data_out <= r_12_2;
		if (write_en==1'b1)
			r_12_2 <= data_in;
	if (addr_selector[12]&addr_selector[3])
		data_out <= r_12_3;
		if (write_en==1'b1)
			r_12_3 <= data_in;
	if (addr_selector[12]&addr_selector[4])
		data_out <= r_12_4;
		if (write_en==1'b1)
			r_12_4 <= data_in;
	if (addr_selector[12]&addr_selector[5])
		data_out <= r_12_5;
		if (write_en==1'b1)
			r_12_5 <= data_in;
	if (addr_selector[12]&addr_selector[6])
		data_out <= r_12_6;
		if (write_en==1'b1)
			r_12_6 <= data_in;
	if (addr_selector[12]&addr_selector[7])
		data_out <= r_12_7;
		if (write_en==1'b1)
			r_12_7 <= data_in;
	if (addr_selector[12]&addr_selector[8])
		data_out <= r_12_8;
		if (write_en==1'b1)
			r_12_8 <= data_in;
	if (addr_selector[12]&addr_selector[9])
		data_out <= r_12_9;
		if (write_en==1'b1)
			r_12_9 <= data_in;
	if (addr_selector[12]&addr_selector[10])
		data_out <= r_12_10;
		if (write_en==1'b1)
			r_12_10 <= data_in;
	if (addr_selector[12]&addr_selector[11])
		data_out <= r_12_11;
		if (write_en==1'b1)
			r_12_11 <= data_in;
	if (addr_selector[12]&addr_selector[12])
		data_out <= r_12_12;
		if (write_en==1'b1)
			r_12_12 <= data_in;
	if (addr_selector[12]&addr_selector[13])
		data_out <= r_12_13;
		if (write_en==1'b1)
			r_12_13 <= data_in;
	if (addr_selector[12]&addr_selector[14])
		data_out <= r_12_14;
		if (write_en==1'b1)
			r_12_14 <= data_in;
	if (addr_selector[12]&addr_selector[15])
		data_out <= r_12_15;
		if (write_en==1'b1)
			r_12_15 <= data_in;
	if (addr_selector[12]&addr_selector[16])
		data_out <= r_12_16;
		if (write_en==1'b1)
			r_12_16 <= data_in;
	if (addr_selector[12]&addr_selector[17])
		data_out <= r_12_17;
		if (write_en==1'b1)
			r_12_17 <= data_in;
	if (addr_selector[12]&addr_selector[18])
		data_out <= r_12_18;
		if (write_en==1'b1)
			r_12_18 <= data_in;
	if (addr_selector[12]&addr_selector[19])
		data_out <= r_12_19;
		if (write_en==1'b1)
			r_12_19 <= data_in;
	if (addr_selector[12]&addr_selector[20])
		data_out <= r_12_20;
		if (write_en==1'b1)
			r_12_20 <= data_in;
	if (addr_selector[12]&addr_selector[21])
		data_out <= r_12_21;
		if (write_en==1'b1)
			r_12_21 <= data_in;
	if (addr_selector[12]&addr_selector[22])
		data_out <= r_12_22;
		if (write_en==1'b1)
			r_12_22 <= data_in;
	if (addr_selector[12]&addr_selector[23])
		data_out <= r_12_23;
		if (write_en==1'b1)
			r_12_23 <= data_in;
	if (addr_selector[12]&addr_selector[24])
		data_out <= r_12_24;
		if (write_en==1'b1)
			r_12_24 <= data_in;
	if (addr_selector[12]&addr_selector[25])
		data_out <= r_12_25;
		if (write_en==1'b1)
			r_12_25 <= data_in;
	if (addr_selector[12]&addr_selector[26])
		data_out <= r_12_26;
		if (write_en==1'b1)
			r_12_26 <= data_in;
	if (addr_selector[12]&addr_selector[27])
		data_out <= r_12_27;
		if (write_en==1'b1)
			r_12_27 <= data_in;
	if (addr_selector[12]&addr_selector[28])
		data_out <= r_12_28;
		if (write_en==1'b1)
			r_12_28 <= data_in;
	if (addr_selector[12]&addr_selector[29])
		data_out <= r_12_29;
		if (write_en==1'b1)
			r_12_29 <= data_in;
	if (addr_selector[12]&addr_selector[30])
		data_out <= r_12_30;
		if (write_en==1'b1)
			r_12_30 <= data_in;
	if (addr_selector[12]&addr_selector[31])
		data_out <= r_12_31;
		if (write_en==1'b1)
			r_12_31 <= data_in;
	if (addr_selector[12]&addr_selector[32])
		data_out <= r_12_32;
		if (write_en==1'b1)
			r_12_32 <= data_in;
	if (addr_selector[12]&addr_selector[33])
		data_out <= r_12_33;
		if (write_en==1'b1)
			r_12_33 <= data_in;
	if (addr_selector[12]&addr_selector[34])
		data_out <= r_12_34;
		if (write_en==1'b1)
			r_12_34 <= data_in;
	if (addr_selector[12]&addr_selector[35])
		data_out <= r_12_35;
		if (write_en==1'b1)
			r_12_35 <= data_in;
	if (addr_selector[12]&addr_selector[36])
		data_out <= r_12_36;
		if (write_en==1'b1)
			r_12_36 <= data_in;
	if (addr_selector[12]&addr_selector[37])
		data_out <= r_12_37;
		if (write_en==1'b1)
			r_12_37 <= data_in;
	if (addr_selector[12]&addr_selector[38])
		data_out <= r_12_38;
		if (write_en==1'b1)
			r_12_38 <= data_in;
	if (addr_selector[12]&addr_selector[39])
		data_out <= r_12_39;
		if (write_en==1'b1)
			r_12_39 <= data_in;
	if (addr_selector[12]&addr_selector[40])
		data_out <= r_12_40;
		if (write_en==1'b1)
			r_12_40 <= data_in;
	if (addr_selector[12]&addr_selector[41])
		data_out <= r_12_41;
		if (write_en==1'b1)
			r_12_41 <= data_in;
	if (addr_selector[12]&addr_selector[42])
		data_out <= r_12_42;
		if (write_en==1'b1)
			r_12_42 <= data_in;
	if (addr_selector[12]&addr_selector[43])
		data_out <= r_12_43;
		if (write_en==1'b1)
			r_12_43 <= data_in;
	if (addr_selector[12]&addr_selector[44])
		data_out <= r_12_44;
		if (write_en==1'b1)
			r_12_44 <= data_in;
	if (addr_selector[12]&addr_selector[45])
		data_out <= r_12_45;
		if (write_en==1'b1)
			r_12_45 <= data_in;
	if (addr_selector[12]&addr_selector[46])
		data_out <= r_12_46;
		if (write_en==1'b1)
			r_12_46 <= data_in;
	if (addr_selector[12]&addr_selector[47])
		data_out <= r_12_47;
		if (write_en==1'b1)
			r_12_47 <= data_in;
	if (addr_selector[12]&addr_selector[48])
		data_out <= r_12_48;
		if (write_en==1'b1)
			r_12_48 <= data_in;
	if (addr_selector[12]&addr_selector[49])
		data_out <= r_12_49;
		if (write_en==1'b1)
			r_12_49 <= data_in;
	if (addr_selector[12]&addr_selector[50])
		data_out <= r_12_50;
		if (write_en==1'b1)
			r_12_50 <= data_in;
	if (addr_selector[12]&addr_selector[51])
		data_out <= r_12_51;
		if (write_en==1'b1)
			r_12_51 <= data_in;
	if (addr_selector[12]&addr_selector[52])
		data_out <= r_12_52;
		if (write_en==1'b1)
			r_12_52 <= data_in;
	if (addr_selector[12]&addr_selector[53])
		data_out <= r_12_53;
		if (write_en==1'b1)
			r_12_53 <= data_in;
	if (addr_selector[12]&addr_selector[54])
		data_out <= r_12_54;
		if (write_en==1'b1)
			r_12_54 <= data_in;
	if (addr_selector[12]&addr_selector[55])
		data_out <= r_12_55;
		if (write_en==1'b1)
			r_12_55 <= data_in;
	if (addr_selector[12]&addr_selector[56])
		data_out <= r_12_56;
		if (write_en==1'b1)
			r_12_56 <= data_in;
	if (addr_selector[12]&addr_selector[57])
		data_out <= r_12_57;
		if (write_en==1'b1)
			r_12_57 <= data_in;
	if (addr_selector[12]&addr_selector[58])
		data_out <= r_12_58;
		if (write_en==1'b1)
			r_12_58 <= data_in;
	if (addr_selector[12]&addr_selector[59])
		data_out <= r_12_59;
		if (write_en==1'b1)
			r_12_59 <= data_in;
	if (addr_selector[12]&addr_selector[60])
		data_out <= r_12_60;
		if (write_en==1'b1)
			r_12_60 <= data_in;
	if (addr_selector[12]&addr_selector[61])
		data_out <= r_12_61;
		if (write_en==1'b1)
			r_12_61 <= data_in;
	if (addr_selector[12]&addr_selector[62])
		data_out <= r_12_62;
		if (write_en==1'b1)
			r_12_62 <= data_in;
	if (addr_selector[12]&addr_selector[63])
		data_out <= r_12_63;
		if (write_en==1'b1)
			r_12_63 <= data_in;
	if (addr_selector[13]&addr_selector[0])
		data_out <= r_13_0;
		if (write_en==1'b1)
			r_13_0 <= data_in;
	if (addr_selector[13]&addr_selector[1])
		data_out <= r_13_1;
		if (write_en==1'b1)
			r_13_1 <= data_in;
	if (addr_selector[13]&addr_selector[2])
		data_out <= r_13_2;
		if (write_en==1'b1)
			r_13_2 <= data_in;
	if (addr_selector[13]&addr_selector[3])
		data_out <= r_13_3;
		if (write_en==1'b1)
			r_13_3 <= data_in;
	if (addr_selector[13]&addr_selector[4])
		data_out <= r_13_4;
		if (write_en==1'b1)
			r_13_4 <= data_in;
	if (addr_selector[13]&addr_selector[5])
		data_out <= r_13_5;
		if (write_en==1'b1)
			r_13_5 <= data_in;
	if (addr_selector[13]&addr_selector[6])
		data_out <= r_13_6;
		if (write_en==1'b1)
			r_13_6 <= data_in;
	if (addr_selector[13]&addr_selector[7])
		data_out <= r_13_7;
		if (write_en==1'b1)
			r_13_7 <= data_in;
	if (addr_selector[13]&addr_selector[8])
		data_out <= r_13_8;
		if (write_en==1'b1)
			r_13_8 <= data_in;
	if (addr_selector[13]&addr_selector[9])
		data_out <= r_13_9;
		if (write_en==1'b1)
			r_13_9 <= data_in;
	if (addr_selector[13]&addr_selector[10])
		data_out <= r_13_10;
		if (write_en==1'b1)
			r_13_10 <= data_in;
	if (addr_selector[13]&addr_selector[11])
		data_out <= r_13_11;
		if (write_en==1'b1)
			r_13_11 <= data_in;
	if (addr_selector[13]&addr_selector[12])
		data_out <= r_13_12;
		if (write_en==1'b1)
			r_13_12 <= data_in;
	if (addr_selector[13]&addr_selector[13])
		data_out <= r_13_13;
		if (write_en==1'b1)
			r_13_13 <= data_in;
	if (addr_selector[13]&addr_selector[14])
		data_out <= r_13_14;
		if (write_en==1'b1)
			r_13_14 <= data_in;
	if (addr_selector[13]&addr_selector[15])
		data_out <= r_13_15;
		if (write_en==1'b1)
			r_13_15 <= data_in;
	if (addr_selector[13]&addr_selector[16])
		data_out <= r_13_16;
		if (write_en==1'b1)
			r_13_16 <= data_in;
	if (addr_selector[13]&addr_selector[17])
		data_out <= r_13_17;
		if (write_en==1'b1)
			r_13_17 <= data_in;
	if (addr_selector[13]&addr_selector[18])
		data_out <= r_13_18;
		if (write_en==1'b1)
			r_13_18 <= data_in;
	if (addr_selector[13]&addr_selector[19])
		data_out <= r_13_19;
		if (write_en==1'b1)
			r_13_19 <= data_in;
	if (addr_selector[13]&addr_selector[20])
		data_out <= r_13_20;
		if (write_en==1'b1)
			r_13_20 <= data_in;
	if (addr_selector[13]&addr_selector[21])
		data_out <= r_13_21;
		if (write_en==1'b1)
			r_13_21 <= data_in;
	if (addr_selector[13]&addr_selector[22])
		data_out <= r_13_22;
		if (write_en==1'b1)
			r_13_22 <= data_in;
	if (addr_selector[13]&addr_selector[23])
		data_out <= r_13_23;
		if (write_en==1'b1)
			r_13_23 <= data_in;
	if (addr_selector[13]&addr_selector[24])
		data_out <= r_13_24;
		if (write_en==1'b1)
			r_13_24 <= data_in;
	if (addr_selector[13]&addr_selector[25])
		data_out <= r_13_25;
		if (write_en==1'b1)
			r_13_25 <= data_in;
	if (addr_selector[13]&addr_selector[26])
		data_out <= r_13_26;
		if (write_en==1'b1)
			r_13_26 <= data_in;
	if (addr_selector[13]&addr_selector[27])
		data_out <= r_13_27;
		if (write_en==1'b1)
			r_13_27 <= data_in;
	if (addr_selector[13]&addr_selector[28])
		data_out <= r_13_28;
		if (write_en==1'b1)
			r_13_28 <= data_in;
	if (addr_selector[13]&addr_selector[29])
		data_out <= r_13_29;
		if (write_en==1'b1)
			r_13_29 <= data_in;
	if (addr_selector[13]&addr_selector[30])
		data_out <= r_13_30;
		if (write_en==1'b1)
			r_13_30 <= data_in;
	if (addr_selector[13]&addr_selector[31])
		data_out <= r_13_31;
		if (write_en==1'b1)
			r_13_31 <= data_in;
	if (addr_selector[13]&addr_selector[32])
		data_out <= r_13_32;
		if (write_en==1'b1)
			r_13_32 <= data_in;
	if (addr_selector[13]&addr_selector[33])
		data_out <= r_13_33;
		if (write_en==1'b1)
			r_13_33 <= data_in;
	if (addr_selector[13]&addr_selector[34])
		data_out <= r_13_34;
		if (write_en==1'b1)
			r_13_34 <= data_in;
	if (addr_selector[13]&addr_selector[35])
		data_out <= r_13_35;
		if (write_en==1'b1)
			r_13_35 <= data_in;
	if (addr_selector[13]&addr_selector[36])
		data_out <= r_13_36;
		if (write_en==1'b1)
			r_13_36 <= data_in;
	if (addr_selector[13]&addr_selector[37])
		data_out <= r_13_37;
		if (write_en==1'b1)
			r_13_37 <= data_in;
	if (addr_selector[13]&addr_selector[38])
		data_out <= r_13_38;
		if (write_en==1'b1)
			r_13_38 <= data_in;
	if (addr_selector[13]&addr_selector[39])
		data_out <= r_13_39;
		if (write_en==1'b1)
			r_13_39 <= data_in;
	if (addr_selector[13]&addr_selector[40])
		data_out <= r_13_40;
		if (write_en==1'b1)
			r_13_40 <= data_in;
	if (addr_selector[13]&addr_selector[41])
		data_out <= r_13_41;
		if (write_en==1'b1)
			r_13_41 <= data_in;
	if (addr_selector[13]&addr_selector[42])
		data_out <= r_13_42;
		if (write_en==1'b1)
			r_13_42 <= data_in;
	if (addr_selector[13]&addr_selector[43])
		data_out <= r_13_43;
		if (write_en==1'b1)
			r_13_43 <= data_in;
	if (addr_selector[13]&addr_selector[44])
		data_out <= r_13_44;
		if (write_en==1'b1)
			r_13_44 <= data_in;
	if (addr_selector[13]&addr_selector[45])
		data_out <= r_13_45;
		if (write_en==1'b1)
			r_13_45 <= data_in;
	if (addr_selector[13]&addr_selector[46])
		data_out <= r_13_46;
		if (write_en==1'b1)
			r_13_46 <= data_in;
	if (addr_selector[13]&addr_selector[47])
		data_out <= r_13_47;
		if (write_en==1'b1)
			r_13_47 <= data_in;
	if (addr_selector[13]&addr_selector[48])
		data_out <= r_13_48;
		if (write_en==1'b1)
			r_13_48 <= data_in;
	if (addr_selector[13]&addr_selector[49])
		data_out <= r_13_49;
		if (write_en==1'b1)
			r_13_49 <= data_in;
	if (addr_selector[13]&addr_selector[50])
		data_out <= r_13_50;
		if (write_en==1'b1)
			r_13_50 <= data_in;
	if (addr_selector[13]&addr_selector[51])
		data_out <= r_13_51;
		if (write_en==1'b1)
			r_13_51 <= data_in;
	if (addr_selector[13]&addr_selector[52])
		data_out <= r_13_52;
		if (write_en==1'b1)
			r_13_52 <= data_in;
	if (addr_selector[13]&addr_selector[53])
		data_out <= r_13_53;
		if (write_en==1'b1)
			r_13_53 <= data_in;
	if (addr_selector[13]&addr_selector[54])
		data_out <= r_13_54;
		if (write_en==1'b1)
			r_13_54 <= data_in;
	if (addr_selector[13]&addr_selector[55])
		data_out <= r_13_55;
		if (write_en==1'b1)
			r_13_55 <= data_in;
	if (addr_selector[13]&addr_selector[56])
		data_out <= r_13_56;
		if (write_en==1'b1)
			r_13_56 <= data_in;
	if (addr_selector[13]&addr_selector[57])
		data_out <= r_13_57;
		if (write_en==1'b1)
			r_13_57 <= data_in;
	if (addr_selector[13]&addr_selector[58])
		data_out <= r_13_58;
		if (write_en==1'b1)
			r_13_58 <= data_in;
	if (addr_selector[13]&addr_selector[59])
		data_out <= r_13_59;
		if (write_en==1'b1)
			r_13_59 <= data_in;
	if (addr_selector[13]&addr_selector[60])
		data_out <= r_13_60;
		if (write_en==1'b1)
			r_13_60 <= data_in;
	if (addr_selector[13]&addr_selector[61])
		data_out <= r_13_61;
		if (write_en==1'b1)
			r_13_61 <= data_in;
	if (addr_selector[13]&addr_selector[62])
		data_out <= r_13_62;
		if (write_en==1'b1)
			r_13_62 <= data_in;
	if (addr_selector[13]&addr_selector[63])
		data_out <= r_13_63;
		if (write_en==1'b1)
			r_13_63 <= data_in;
	if (addr_selector[14]&addr_selector[0])
		data_out <= r_14_0;
		if (write_en==1'b1)
			r_14_0 <= data_in;
	if (addr_selector[14]&addr_selector[1])
		data_out <= r_14_1;
		if (write_en==1'b1)
			r_14_1 <= data_in;
	if (addr_selector[14]&addr_selector[2])
		data_out <= r_14_2;
		if (write_en==1'b1)
			r_14_2 <= data_in;
	if (addr_selector[14]&addr_selector[3])
		data_out <= r_14_3;
		if (write_en==1'b1)
			r_14_3 <= data_in;
	if (addr_selector[14]&addr_selector[4])
		data_out <= r_14_4;
		if (write_en==1'b1)
			r_14_4 <= data_in;
	if (addr_selector[14]&addr_selector[5])
		data_out <= r_14_5;
		if (write_en==1'b1)
			r_14_5 <= data_in;
	if (addr_selector[14]&addr_selector[6])
		data_out <= r_14_6;
		if (write_en==1'b1)
			r_14_6 <= data_in;
	if (addr_selector[14]&addr_selector[7])
		data_out <= r_14_7;
		if (write_en==1'b1)
			r_14_7 <= data_in;
	if (addr_selector[14]&addr_selector[8])
		data_out <= r_14_8;
		if (write_en==1'b1)
			r_14_8 <= data_in;
	if (addr_selector[14]&addr_selector[9])
		data_out <= r_14_9;
		if (write_en==1'b1)
			r_14_9 <= data_in;
	if (addr_selector[14]&addr_selector[10])
		data_out <= r_14_10;
		if (write_en==1'b1)
			r_14_10 <= data_in;
	if (addr_selector[14]&addr_selector[11])
		data_out <= r_14_11;
		if (write_en==1'b1)
			r_14_11 <= data_in;
	if (addr_selector[14]&addr_selector[12])
		data_out <= r_14_12;
		if (write_en==1'b1)
			r_14_12 <= data_in;
	if (addr_selector[14]&addr_selector[13])
		data_out <= r_14_13;
		if (write_en==1'b1)
			r_14_13 <= data_in;
	if (addr_selector[14]&addr_selector[14])
		data_out <= r_14_14;
		if (write_en==1'b1)
			r_14_14 <= data_in;
	if (addr_selector[14]&addr_selector[15])
		data_out <= r_14_15;
		if (write_en==1'b1)
			r_14_15 <= data_in;
	if (addr_selector[14]&addr_selector[16])
		data_out <= r_14_16;
		if (write_en==1'b1)
			r_14_16 <= data_in;
	if (addr_selector[14]&addr_selector[17])
		data_out <= r_14_17;
		if (write_en==1'b1)
			r_14_17 <= data_in;
	if (addr_selector[14]&addr_selector[18])
		data_out <= r_14_18;
		if (write_en==1'b1)
			r_14_18 <= data_in;
	if (addr_selector[14]&addr_selector[19])
		data_out <= r_14_19;
		if (write_en==1'b1)
			r_14_19 <= data_in;
	if (addr_selector[14]&addr_selector[20])
		data_out <= r_14_20;
		if (write_en==1'b1)
			r_14_20 <= data_in;
	if (addr_selector[14]&addr_selector[21])
		data_out <= r_14_21;
		if (write_en==1'b1)
			r_14_21 <= data_in;
	if (addr_selector[14]&addr_selector[22])
		data_out <= r_14_22;
		if (write_en==1'b1)
			r_14_22 <= data_in;
	if (addr_selector[14]&addr_selector[23])
		data_out <= r_14_23;
		if (write_en==1'b1)
			r_14_23 <= data_in;
	if (addr_selector[14]&addr_selector[24])
		data_out <= r_14_24;
		if (write_en==1'b1)
			r_14_24 <= data_in;
	if (addr_selector[14]&addr_selector[25])
		data_out <= r_14_25;
		if (write_en==1'b1)
			r_14_25 <= data_in;
	if (addr_selector[14]&addr_selector[26])
		data_out <= r_14_26;
		if (write_en==1'b1)
			r_14_26 <= data_in;
	if (addr_selector[14]&addr_selector[27])
		data_out <= r_14_27;
		if (write_en==1'b1)
			r_14_27 <= data_in;
	if (addr_selector[14]&addr_selector[28])
		data_out <= r_14_28;
		if (write_en==1'b1)
			r_14_28 <= data_in;
	if (addr_selector[14]&addr_selector[29])
		data_out <= r_14_29;
		if (write_en==1'b1)
			r_14_29 <= data_in;
	if (addr_selector[14]&addr_selector[30])
		data_out <= r_14_30;
		if (write_en==1'b1)
			r_14_30 <= data_in;
	if (addr_selector[14]&addr_selector[31])
		data_out <= r_14_31;
		if (write_en==1'b1)
			r_14_31 <= data_in;
	if (addr_selector[14]&addr_selector[32])
		data_out <= r_14_32;
		if (write_en==1'b1)
			r_14_32 <= data_in;
	if (addr_selector[14]&addr_selector[33])
		data_out <= r_14_33;
		if (write_en==1'b1)
			r_14_33 <= data_in;
	if (addr_selector[14]&addr_selector[34])
		data_out <= r_14_34;
		if (write_en==1'b1)
			r_14_34 <= data_in;
	if (addr_selector[14]&addr_selector[35])
		data_out <= r_14_35;
		if (write_en==1'b1)
			r_14_35 <= data_in;
	if (addr_selector[14]&addr_selector[36])
		data_out <= r_14_36;
		if (write_en==1'b1)
			r_14_36 <= data_in;
	if (addr_selector[14]&addr_selector[37])
		data_out <= r_14_37;
		if (write_en==1'b1)
			r_14_37 <= data_in;
	if (addr_selector[14]&addr_selector[38])
		data_out <= r_14_38;
		if (write_en==1'b1)
			r_14_38 <= data_in;
	if (addr_selector[14]&addr_selector[39])
		data_out <= r_14_39;
		if (write_en==1'b1)
			r_14_39 <= data_in;
	if (addr_selector[14]&addr_selector[40])
		data_out <= r_14_40;
		if (write_en==1'b1)
			r_14_40 <= data_in;
	if (addr_selector[14]&addr_selector[41])
		data_out <= r_14_41;
		if (write_en==1'b1)
			r_14_41 <= data_in;
	if (addr_selector[14]&addr_selector[42])
		data_out <= r_14_42;
		if (write_en==1'b1)
			r_14_42 <= data_in;
	if (addr_selector[14]&addr_selector[43])
		data_out <= r_14_43;
		if (write_en==1'b1)
			r_14_43 <= data_in;
	if (addr_selector[14]&addr_selector[44])
		data_out <= r_14_44;
		if (write_en==1'b1)
			r_14_44 <= data_in;
	if (addr_selector[14]&addr_selector[45])
		data_out <= r_14_45;
		if (write_en==1'b1)
			r_14_45 <= data_in;
	if (addr_selector[14]&addr_selector[46])
		data_out <= r_14_46;
		if (write_en==1'b1)
			r_14_46 <= data_in;
	if (addr_selector[14]&addr_selector[47])
		data_out <= r_14_47;
		if (write_en==1'b1)
			r_14_47 <= data_in;
	if (addr_selector[14]&addr_selector[48])
		data_out <= r_14_48;
		if (write_en==1'b1)
			r_14_48 <= data_in;
	if (addr_selector[14]&addr_selector[49])
		data_out <= r_14_49;
		if (write_en==1'b1)
			r_14_49 <= data_in;
	if (addr_selector[14]&addr_selector[50])
		data_out <= r_14_50;
		if (write_en==1'b1)
			r_14_50 <= data_in;
	if (addr_selector[14]&addr_selector[51])
		data_out <= r_14_51;
		if (write_en==1'b1)
			r_14_51 <= data_in;
	if (addr_selector[14]&addr_selector[52])
		data_out <= r_14_52;
		if (write_en==1'b1)
			r_14_52 <= data_in;
	if (addr_selector[14]&addr_selector[53])
		data_out <= r_14_53;
		if (write_en==1'b1)
			r_14_53 <= data_in;
	if (addr_selector[14]&addr_selector[54])
		data_out <= r_14_54;
		if (write_en==1'b1)
			r_14_54 <= data_in;
	if (addr_selector[14]&addr_selector[55])
		data_out <= r_14_55;
		if (write_en==1'b1)
			r_14_55 <= data_in;
	if (addr_selector[14]&addr_selector[56])
		data_out <= r_14_56;
		if (write_en==1'b1)
			r_14_56 <= data_in;
	if (addr_selector[14]&addr_selector[57])
		data_out <= r_14_57;
		if (write_en==1'b1)
			r_14_57 <= data_in;
	if (addr_selector[14]&addr_selector[58])
		data_out <= r_14_58;
		if (write_en==1'b1)
			r_14_58 <= data_in;
	if (addr_selector[14]&addr_selector[59])
		data_out <= r_14_59;
		if (write_en==1'b1)
			r_14_59 <= data_in;
	if (addr_selector[14]&addr_selector[60])
		data_out <= r_14_60;
		if (write_en==1'b1)
			r_14_60 <= data_in;
	if (addr_selector[14]&addr_selector[61])
		data_out <= r_14_61;
		if (write_en==1'b1)
			r_14_61 <= data_in;
	if (addr_selector[14]&addr_selector[62])
		data_out <= r_14_62;
		if (write_en==1'b1)
			r_14_62 <= data_in;
	if (addr_selector[14]&addr_selector[63])
		data_out <= r_14_63;
		if (write_en==1'b1)
			r_14_63 <= data_in;
	if (addr_selector[15]&addr_selector[0])
		data_out <= r_15_0;
		if (write_en==1'b1)
			r_15_0 <= data_in;
	if (addr_selector[15]&addr_selector[1])
		data_out <= r_15_1;
		if (write_en==1'b1)
			r_15_1 <= data_in;
	if (addr_selector[15]&addr_selector[2])
		data_out <= r_15_2;
		if (write_en==1'b1)
			r_15_2 <= data_in;
	if (addr_selector[15]&addr_selector[3])
		data_out <= r_15_3;
		if (write_en==1'b1)
			r_15_3 <= data_in;
	if (addr_selector[15]&addr_selector[4])
		data_out <= r_15_4;
		if (write_en==1'b1)
			r_15_4 <= data_in;
	if (addr_selector[15]&addr_selector[5])
		data_out <= r_15_5;
		if (write_en==1'b1)
			r_15_5 <= data_in;
	if (addr_selector[15]&addr_selector[6])
		data_out <= r_15_6;
		if (write_en==1'b1)
			r_15_6 <= data_in;
	if (addr_selector[15]&addr_selector[7])
		data_out <= r_15_7;
		if (write_en==1'b1)
			r_15_7 <= data_in;
	if (addr_selector[15]&addr_selector[8])
		data_out <= r_15_8;
		if (write_en==1'b1)
			r_15_8 <= data_in;
	if (addr_selector[15]&addr_selector[9])
		data_out <= r_15_9;
		if (write_en==1'b1)
			r_15_9 <= data_in;
	if (addr_selector[15]&addr_selector[10])
		data_out <= r_15_10;
		if (write_en==1'b1)
			r_15_10 <= data_in;
	if (addr_selector[15]&addr_selector[11])
		data_out <= r_15_11;
		if (write_en==1'b1)
			r_15_11 <= data_in;
	if (addr_selector[15]&addr_selector[12])
		data_out <= r_15_12;
		if (write_en==1'b1)
			r_15_12 <= data_in;
	if (addr_selector[15]&addr_selector[13])
		data_out <= r_15_13;
		if (write_en==1'b1)
			r_15_13 <= data_in;
	if (addr_selector[15]&addr_selector[14])
		data_out <= r_15_14;
		if (write_en==1'b1)
			r_15_14 <= data_in;
	if (addr_selector[15]&addr_selector[15])
		data_out <= r_15_15;
		if (write_en==1'b1)
			r_15_15 <= data_in;
	if (addr_selector[15]&addr_selector[16])
		data_out <= r_15_16;
		if (write_en==1'b1)
			r_15_16 <= data_in;
	if (addr_selector[15]&addr_selector[17])
		data_out <= r_15_17;
		if (write_en==1'b1)
			r_15_17 <= data_in;
	if (addr_selector[15]&addr_selector[18])
		data_out <= r_15_18;
		if (write_en==1'b1)
			r_15_18 <= data_in;
	if (addr_selector[15]&addr_selector[19])
		data_out <= r_15_19;
		if (write_en==1'b1)
			r_15_19 <= data_in;
	if (addr_selector[15]&addr_selector[20])
		data_out <= r_15_20;
		if (write_en==1'b1)
			r_15_20 <= data_in;
	if (addr_selector[15]&addr_selector[21])
		data_out <= r_15_21;
		if (write_en==1'b1)
			r_15_21 <= data_in;
	if (addr_selector[15]&addr_selector[22])
		data_out <= r_15_22;
		if (write_en==1'b1)
			r_15_22 <= data_in;
	if (addr_selector[15]&addr_selector[23])
		data_out <= r_15_23;
		if (write_en==1'b1)
			r_15_23 <= data_in;
	if (addr_selector[15]&addr_selector[24])
		data_out <= r_15_24;
		if (write_en==1'b1)
			r_15_24 <= data_in;
	if (addr_selector[15]&addr_selector[25])
		data_out <= r_15_25;
		if (write_en==1'b1)
			r_15_25 <= data_in;
	if (addr_selector[15]&addr_selector[26])
		data_out <= r_15_26;
		if (write_en==1'b1)
			r_15_26 <= data_in;
	if (addr_selector[15]&addr_selector[27])
		data_out <= r_15_27;
		if (write_en==1'b1)
			r_15_27 <= data_in;
	if (addr_selector[15]&addr_selector[28])
		data_out <= r_15_28;
		if (write_en==1'b1)
			r_15_28 <= data_in;
	if (addr_selector[15]&addr_selector[29])
		data_out <= r_15_29;
		if (write_en==1'b1)
			r_15_29 <= data_in;
	if (addr_selector[15]&addr_selector[30])
		data_out <= r_15_30;
		if (write_en==1'b1)
			r_15_30 <= data_in;
	if (addr_selector[15]&addr_selector[31])
		data_out <= r_15_31;
		if (write_en==1'b1)
			r_15_31 <= data_in;
	if (addr_selector[15]&addr_selector[32])
		data_out <= r_15_32;
		if (write_en==1'b1)
			r_15_32 <= data_in;
	if (addr_selector[15]&addr_selector[33])
		data_out <= r_15_33;
		if (write_en==1'b1)
			r_15_33 <= data_in;
	if (addr_selector[15]&addr_selector[34])
		data_out <= r_15_34;
		if (write_en==1'b1)
			r_15_34 <= data_in;
	if (addr_selector[15]&addr_selector[35])
		data_out <= r_15_35;
		if (write_en==1'b1)
			r_15_35 <= data_in;
	if (addr_selector[15]&addr_selector[36])
		data_out <= r_15_36;
		if (write_en==1'b1)
			r_15_36 <= data_in;
	if (addr_selector[15]&addr_selector[37])
		data_out <= r_15_37;
		if (write_en==1'b1)
			r_15_37 <= data_in;
	if (addr_selector[15]&addr_selector[38])
		data_out <= r_15_38;
		if (write_en==1'b1)
			r_15_38 <= data_in;
	if (addr_selector[15]&addr_selector[39])
		data_out <= r_15_39;
		if (write_en==1'b1)
			r_15_39 <= data_in;
	if (addr_selector[15]&addr_selector[40])
		data_out <= r_15_40;
		if (write_en==1'b1)
			r_15_40 <= data_in;
	if (addr_selector[15]&addr_selector[41])
		data_out <= r_15_41;
		if (write_en==1'b1)
			r_15_41 <= data_in;
	if (addr_selector[15]&addr_selector[42])
		data_out <= r_15_42;
		if (write_en==1'b1)
			r_15_42 <= data_in;
	if (addr_selector[15]&addr_selector[43])
		data_out <= r_15_43;
		if (write_en==1'b1)
			r_15_43 <= data_in;
	if (addr_selector[15]&addr_selector[44])
		data_out <= r_15_44;
		if (write_en==1'b1)
			r_15_44 <= data_in;
	if (addr_selector[15]&addr_selector[45])
		data_out <= r_15_45;
		if (write_en==1'b1)
			r_15_45 <= data_in;
	if (addr_selector[15]&addr_selector[46])
		data_out <= r_15_46;
		if (write_en==1'b1)
			r_15_46 <= data_in;
	if (addr_selector[15]&addr_selector[47])
		data_out <= r_15_47;
		if (write_en==1'b1)
			r_15_47 <= data_in;
	if (addr_selector[15]&addr_selector[48])
		data_out <= r_15_48;
		if (write_en==1'b1)
			r_15_48 <= data_in;
	if (addr_selector[15]&addr_selector[49])
		data_out <= r_15_49;
		if (write_en==1'b1)
			r_15_49 <= data_in;
	if (addr_selector[15]&addr_selector[50])
		data_out <= r_15_50;
		if (write_en==1'b1)
			r_15_50 <= data_in;
	if (addr_selector[15]&addr_selector[51])
		data_out <= r_15_51;
		if (write_en==1'b1)
			r_15_51 <= data_in;
	if (addr_selector[15]&addr_selector[52])
		data_out <= r_15_52;
		if (write_en==1'b1)
			r_15_52 <= data_in;
	if (addr_selector[15]&addr_selector[53])
		data_out <= r_15_53;
		if (write_en==1'b1)
			r_15_53 <= data_in;
	if (addr_selector[15]&addr_selector[54])
		data_out <= r_15_54;
		if (write_en==1'b1)
			r_15_54 <= data_in;
	if (addr_selector[15]&addr_selector[55])
		data_out <= r_15_55;
		if (write_en==1'b1)
			r_15_55 <= data_in;
	if (addr_selector[15]&addr_selector[56])
		data_out <= r_15_56;
		if (write_en==1'b1)
			r_15_56 <= data_in;
	if (addr_selector[15]&addr_selector[57])
		data_out <= r_15_57;
		if (write_en==1'b1)
			r_15_57 <= data_in;
	if (addr_selector[15]&addr_selector[58])
		data_out <= r_15_58;
		if (write_en==1'b1)
			r_15_58 <= data_in;
	if (addr_selector[15]&addr_selector[59])
		data_out <= r_15_59;
		if (write_en==1'b1)
			r_15_59 <= data_in;
	if (addr_selector[15]&addr_selector[60])
		data_out <= r_15_60;
		if (write_en==1'b1)
			r_15_60 <= data_in;
	if (addr_selector[15]&addr_selector[61])
		data_out <= r_15_61;
		if (write_en==1'b1)
			r_15_61 <= data_in;
	if (addr_selector[15]&addr_selector[62])
		data_out <= r_15_62;
		if (write_en==1'b1)
			r_15_62 <= data_in;
	if (addr_selector[15]&addr_selector[63])
		data_out <= r_15_63;
		if (write_en==1'b1)
			r_15_63 <= data_in;
	if (addr_selector[16]&addr_selector[0])
		data_out <= r_16_0;
		if (write_en==1'b1)
			r_16_0 <= data_in;
	if (addr_selector[16]&addr_selector[1])
		data_out <= r_16_1;
		if (write_en==1'b1)
			r_16_1 <= data_in;
	if (addr_selector[16]&addr_selector[2])
		data_out <= r_16_2;
		if (write_en==1'b1)
			r_16_2 <= data_in;
	if (addr_selector[16]&addr_selector[3])
		data_out <= r_16_3;
		if (write_en==1'b1)
			r_16_3 <= data_in;
	if (addr_selector[16]&addr_selector[4])
		data_out <= r_16_4;
		if (write_en==1'b1)
			r_16_4 <= data_in;
	if (addr_selector[16]&addr_selector[5])
		data_out <= r_16_5;
		if (write_en==1'b1)
			r_16_5 <= data_in;
	if (addr_selector[16]&addr_selector[6])
		data_out <= r_16_6;
		if (write_en==1'b1)
			r_16_6 <= data_in;
	if (addr_selector[16]&addr_selector[7])
		data_out <= r_16_7;
		if (write_en==1'b1)
			r_16_7 <= data_in;
	if (addr_selector[16]&addr_selector[8])
		data_out <= r_16_8;
		if (write_en==1'b1)
			r_16_8 <= data_in;
	if (addr_selector[16]&addr_selector[9])
		data_out <= r_16_9;
		if (write_en==1'b1)
			r_16_9 <= data_in;
	if (addr_selector[16]&addr_selector[10])
		data_out <= r_16_10;
		if (write_en==1'b1)
			r_16_10 <= data_in;
	if (addr_selector[16]&addr_selector[11])
		data_out <= r_16_11;
		if (write_en==1'b1)
			r_16_11 <= data_in;
	if (addr_selector[16]&addr_selector[12])
		data_out <= r_16_12;
		if (write_en==1'b1)
			r_16_12 <= data_in;
	if (addr_selector[16]&addr_selector[13])
		data_out <= r_16_13;
		if (write_en==1'b1)
			r_16_13 <= data_in;
	if (addr_selector[16]&addr_selector[14])
		data_out <= r_16_14;
		if (write_en==1'b1)
			r_16_14 <= data_in;
	if (addr_selector[16]&addr_selector[15])
		data_out <= r_16_15;
		if (write_en==1'b1)
			r_16_15 <= data_in;
	if (addr_selector[16]&addr_selector[16])
		data_out <= r_16_16;
		if (write_en==1'b1)
			r_16_16 <= data_in;
	if (addr_selector[16]&addr_selector[17])
		data_out <= r_16_17;
		if (write_en==1'b1)
			r_16_17 <= data_in;
	if (addr_selector[16]&addr_selector[18])
		data_out <= r_16_18;
		if (write_en==1'b1)
			r_16_18 <= data_in;
	if (addr_selector[16]&addr_selector[19])
		data_out <= r_16_19;
		if (write_en==1'b1)
			r_16_19 <= data_in;
	if (addr_selector[16]&addr_selector[20])
		data_out <= r_16_20;
		if (write_en==1'b1)
			r_16_20 <= data_in;
	if (addr_selector[16]&addr_selector[21])
		data_out <= r_16_21;
		if (write_en==1'b1)
			r_16_21 <= data_in;
	if (addr_selector[16]&addr_selector[22])
		data_out <= r_16_22;
		if (write_en==1'b1)
			r_16_22 <= data_in;
	if (addr_selector[16]&addr_selector[23])
		data_out <= r_16_23;
		if (write_en==1'b1)
			r_16_23 <= data_in;
	if (addr_selector[16]&addr_selector[24])
		data_out <= r_16_24;
		if (write_en==1'b1)
			r_16_24 <= data_in;
	if (addr_selector[16]&addr_selector[25])
		data_out <= r_16_25;
		if (write_en==1'b1)
			r_16_25 <= data_in;
	if (addr_selector[16]&addr_selector[26])
		data_out <= r_16_26;
		if (write_en==1'b1)
			r_16_26 <= data_in;
	if (addr_selector[16]&addr_selector[27])
		data_out <= r_16_27;
		if (write_en==1'b1)
			r_16_27 <= data_in;
	if (addr_selector[16]&addr_selector[28])
		data_out <= r_16_28;
		if (write_en==1'b1)
			r_16_28 <= data_in;
	if (addr_selector[16]&addr_selector[29])
		data_out <= r_16_29;
		if (write_en==1'b1)
			r_16_29 <= data_in;
	if (addr_selector[16]&addr_selector[30])
		data_out <= r_16_30;
		if (write_en==1'b1)
			r_16_30 <= data_in;
	if (addr_selector[16]&addr_selector[31])
		data_out <= r_16_31;
		if (write_en==1'b1)
			r_16_31 <= data_in;
	if (addr_selector[16]&addr_selector[32])
		data_out <= r_16_32;
		if (write_en==1'b1)
			r_16_32 <= data_in;
	if (addr_selector[16]&addr_selector[33])
		data_out <= r_16_33;
		if (write_en==1'b1)
			r_16_33 <= data_in;
	if (addr_selector[16]&addr_selector[34])
		data_out <= r_16_34;
		if (write_en==1'b1)
			r_16_34 <= data_in;
	if (addr_selector[16]&addr_selector[35])
		data_out <= r_16_35;
		if (write_en==1'b1)
			r_16_35 <= data_in;
	if (addr_selector[16]&addr_selector[36])
		data_out <= r_16_36;
		if (write_en==1'b1)
			r_16_36 <= data_in;
	if (addr_selector[16]&addr_selector[37])
		data_out <= r_16_37;
		if (write_en==1'b1)
			r_16_37 <= data_in;
	if (addr_selector[16]&addr_selector[38])
		data_out <= r_16_38;
		if (write_en==1'b1)
			r_16_38 <= data_in;
	if (addr_selector[16]&addr_selector[39])
		data_out <= r_16_39;
		if (write_en==1'b1)
			r_16_39 <= data_in;
	if (addr_selector[16]&addr_selector[40])
		data_out <= r_16_40;
		if (write_en==1'b1)
			r_16_40 <= data_in;
	if (addr_selector[16]&addr_selector[41])
		data_out <= r_16_41;
		if (write_en==1'b1)
			r_16_41 <= data_in;
	if (addr_selector[16]&addr_selector[42])
		data_out <= r_16_42;
		if (write_en==1'b1)
			r_16_42 <= data_in;
	if (addr_selector[16]&addr_selector[43])
		data_out <= r_16_43;
		if (write_en==1'b1)
			r_16_43 <= data_in;
	if (addr_selector[16]&addr_selector[44])
		data_out <= r_16_44;
		if (write_en==1'b1)
			r_16_44 <= data_in;
	if (addr_selector[16]&addr_selector[45])
		data_out <= r_16_45;
		if (write_en==1'b1)
			r_16_45 <= data_in;
	if (addr_selector[16]&addr_selector[46])
		data_out <= r_16_46;
		if (write_en==1'b1)
			r_16_46 <= data_in;
	if (addr_selector[16]&addr_selector[47])
		data_out <= r_16_47;
		if (write_en==1'b1)
			r_16_47 <= data_in;
	if (addr_selector[16]&addr_selector[48])
		data_out <= r_16_48;
		if (write_en==1'b1)
			r_16_48 <= data_in;
	if (addr_selector[16]&addr_selector[49])
		data_out <= r_16_49;
		if (write_en==1'b1)
			r_16_49 <= data_in;
	if (addr_selector[16]&addr_selector[50])
		data_out <= r_16_50;
		if (write_en==1'b1)
			r_16_50 <= data_in;
	if (addr_selector[16]&addr_selector[51])
		data_out <= r_16_51;
		if (write_en==1'b1)
			r_16_51 <= data_in;
	if (addr_selector[16]&addr_selector[52])
		data_out <= r_16_52;
		if (write_en==1'b1)
			r_16_52 <= data_in;
	if (addr_selector[16]&addr_selector[53])
		data_out <= r_16_53;
		if (write_en==1'b1)
			r_16_53 <= data_in;
	if (addr_selector[16]&addr_selector[54])
		data_out <= r_16_54;
		if (write_en==1'b1)
			r_16_54 <= data_in;
	if (addr_selector[16]&addr_selector[55])
		data_out <= r_16_55;
		if (write_en==1'b1)
			r_16_55 <= data_in;
	if (addr_selector[16]&addr_selector[56])
		data_out <= r_16_56;
		if (write_en==1'b1)
			r_16_56 <= data_in;
	if (addr_selector[16]&addr_selector[57])
		data_out <= r_16_57;
		if (write_en==1'b1)
			r_16_57 <= data_in;
	if (addr_selector[16]&addr_selector[58])
		data_out <= r_16_58;
		if (write_en==1'b1)
			r_16_58 <= data_in;
	if (addr_selector[16]&addr_selector[59])
		data_out <= r_16_59;
		if (write_en==1'b1)
			r_16_59 <= data_in;
	if (addr_selector[16]&addr_selector[60])
		data_out <= r_16_60;
		if (write_en==1'b1)
			r_16_60 <= data_in;
	if (addr_selector[16]&addr_selector[61])
		data_out <= r_16_61;
		if (write_en==1'b1)
			r_16_61 <= data_in;
	if (addr_selector[16]&addr_selector[62])
		data_out <= r_16_62;
		if (write_en==1'b1)
			r_16_62 <= data_in;
	if (addr_selector[16]&addr_selector[63])
		data_out <= r_16_63;
		if (write_en==1'b1)
			r_16_63 <= data_in;
	if (addr_selector[17]&addr_selector[0])
		data_out <= r_17_0;
		if (write_en==1'b1)
			r_17_0 <= data_in;
	if (addr_selector[17]&addr_selector[1])
		data_out <= r_17_1;
		if (write_en==1'b1)
			r_17_1 <= data_in;
	if (addr_selector[17]&addr_selector[2])
		data_out <= r_17_2;
		if (write_en==1'b1)
			r_17_2 <= data_in;
	if (addr_selector[17]&addr_selector[3])
		data_out <= r_17_3;
		if (write_en==1'b1)
			r_17_3 <= data_in;
	if (addr_selector[17]&addr_selector[4])
		data_out <= r_17_4;
		if (write_en==1'b1)
			r_17_4 <= data_in;
	if (addr_selector[17]&addr_selector[5])
		data_out <= r_17_5;
		if (write_en==1'b1)
			r_17_5 <= data_in;
	if (addr_selector[17]&addr_selector[6])
		data_out <= r_17_6;
		if (write_en==1'b1)
			r_17_6 <= data_in;
	if (addr_selector[17]&addr_selector[7])
		data_out <= r_17_7;
		if (write_en==1'b1)
			r_17_7 <= data_in;
	if (addr_selector[17]&addr_selector[8])
		data_out <= r_17_8;
		if (write_en==1'b1)
			r_17_8 <= data_in;
	if (addr_selector[17]&addr_selector[9])
		data_out <= r_17_9;
		if (write_en==1'b1)
			r_17_9 <= data_in;
	if (addr_selector[17]&addr_selector[10])
		data_out <= r_17_10;
		if (write_en==1'b1)
			r_17_10 <= data_in;
	if (addr_selector[17]&addr_selector[11])
		data_out <= r_17_11;
		if (write_en==1'b1)
			r_17_11 <= data_in;
	if (addr_selector[17]&addr_selector[12])
		data_out <= r_17_12;
		if (write_en==1'b1)
			r_17_12 <= data_in;
	if (addr_selector[17]&addr_selector[13])
		data_out <= r_17_13;
		if (write_en==1'b1)
			r_17_13 <= data_in;
	if (addr_selector[17]&addr_selector[14])
		data_out <= r_17_14;
		if (write_en==1'b1)
			r_17_14 <= data_in;
	if (addr_selector[17]&addr_selector[15])
		data_out <= r_17_15;
		if (write_en==1'b1)
			r_17_15 <= data_in;
	if (addr_selector[17]&addr_selector[16])
		data_out <= r_17_16;
		if (write_en==1'b1)
			r_17_16 <= data_in;
	if (addr_selector[17]&addr_selector[17])
		data_out <= r_17_17;
		if (write_en==1'b1)
			r_17_17 <= data_in;
	if (addr_selector[17]&addr_selector[18])
		data_out <= r_17_18;
		if (write_en==1'b1)
			r_17_18 <= data_in;
	if (addr_selector[17]&addr_selector[19])
		data_out <= r_17_19;
		if (write_en==1'b1)
			r_17_19 <= data_in;
	if (addr_selector[17]&addr_selector[20])
		data_out <= r_17_20;
		if (write_en==1'b1)
			r_17_20 <= data_in;
	if (addr_selector[17]&addr_selector[21])
		data_out <= r_17_21;
		if (write_en==1'b1)
			r_17_21 <= data_in;
	if (addr_selector[17]&addr_selector[22])
		data_out <= r_17_22;
		if (write_en==1'b1)
			r_17_22 <= data_in;
	if (addr_selector[17]&addr_selector[23])
		data_out <= r_17_23;
		if (write_en==1'b1)
			r_17_23 <= data_in;
	if (addr_selector[17]&addr_selector[24])
		data_out <= r_17_24;
		if (write_en==1'b1)
			r_17_24 <= data_in;
	if (addr_selector[17]&addr_selector[25])
		data_out <= r_17_25;
		if (write_en==1'b1)
			r_17_25 <= data_in;
	if (addr_selector[17]&addr_selector[26])
		data_out <= r_17_26;
		if (write_en==1'b1)
			r_17_26 <= data_in;
	if (addr_selector[17]&addr_selector[27])
		data_out <= r_17_27;
		if (write_en==1'b1)
			r_17_27 <= data_in;
	if (addr_selector[17]&addr_selector[28])
		data_out <= r_17_28;
		if (write_en==1'b1)
			r_17_28 <= data_in;
	if (addr_selector[17]&addr_selector[29])
		data_out <= r_17_29;
		if (write_en==1'b1)
			r_17_29 <= data_in;
	if (addr_selector[17]&addr_selector[30])
		data_out <= r_17_30;
		if (write_en==1'b1)
			r_17_30 <= data_in;
	if (addr_selector[17]&addr_selector[31])
		data_out <= r_17_31;
		if (write_en==1'b1)
			r_17_31 <= data_in;
	if (addr_selector[17]&addr_selector[32])
		data_out <= r_17_32;
		if (write_en==1'b1)
			r_17_32 <= data_in;
	if (addr_selector[17]&addr_selector[33])
		data_out <= r_17_33;
		if (write_en==1'b1)
			r_17_33 <= data_in;
	if (addr_selector[17]&addr_selector[34])
		data_out <= r_17_34;
		if (write_en==1'b1)
			r_17_34 <= data_in;
	if (addr_selector[17]&addr_selector[35])
		data_out <= r_17_35;
		if (write_en==1'b1)
			r_17_35 <= data_in;
	if (addr_selector[17]&addr_selector[36])
		data_out <= r_17_36;
		if (write_en==1'b1)
			r_17_36 <= data_in;
	if (addr_selector[17]&addr_selector[37])
		data_out <= r_17_37;
		if (write_en==1'b1)
			r_17_37 <= data_in;
	if (addr_selector[17]&addr_selector[38])
		data_out <= r_17_38;
		if (write_en==1'b1)
			r_17_38 <= data_in;
	if (addr_selector[17]&addr_selector[39])
		data_out <= r_17_39;
		if (write_en==1'b1)
			r_17_39 <= data_in;
	if (addr_selector[17]&addr_selector[40])
		data_out <= r_17_40;
		if (write_en==1'b1)
			r_17_40 <= data_in;
	if (addr_selector[17]&addr_selector[41])
		data_out <= r_17_41;
		if (write_en==1'b1)
			r_17_41 <= data_in;
	if (addr_selector[17]&addr_selector[42])
		data_out <= r_17_42;
		if (write_en==1'b1)
			r_17_42 <= data_in;
	if (addr_selector[17]&addr_selector[43])
		data_out <= r_17_43;
		if (write_en==1'b1)
			r_17_43 <= data_in;
	if (addr_selector[17]&addr_selector[44])
		data_out <= r_17_44;
		if (write_en==1'b1)
			r_17_44 <= data_in;
	if (addr_selector[17]&addr_selector[45])
		data_out <= r_17_45;
		if (write_en==1'b1)
			r_17_45 <= data_in;
	if (addr_selector[17]&addr_selector[46])
		data_out <= r_17_46;
		if (write_en==1'b1)
			r_17_46 <= data_in;
	if (addr_selector[17]&addr_selector[47])
		data_out <= r_17_47;
		if (write_en==1'b1)
			r_17_47 <= data_in;
	if (addr_selector[17]&addr_selector[48])
		data_out <= r_17_48;
		if (write_en==1'b1)
			r_17_48 <= data_in;
	if (addr_selector[17]&addr_selector[49])
		data_out <= r_17_49;
		if (write_en==1'b1)
			r_17_49 <= data_in;
	if (addr_selector[17]&addr_selector[50])
		data_out <= r_17_50;
		if (write_en==1'b1)
			r_17_50 <= data_in;
	if (addr_selector[17]&addr_selector[51])
		data_out <= r_17_51;
		if (write_en==1'b1)
			r_17_51 <= data_in;
	if (addr_selector[17]&addr_selector[52])
		data_out <= r_17_52;
		if (write_en==1'b1)
			r_17_52 <= data_in;
	if (addr_selector[17]&addr_selector[53])
		data_out <= r_17_53;
		if (write_en==1'b1)
			r_17_53 <= data_in;
	if (addr_selector[17]&addr_selector[54])
		data_out <= r_17_54;
		if (write_en==1'b1)
			r_17_54 <= data_in;
	if (addr_selector[17]&addr_selector[55])
		data_out <= r_17_55;
		if (write_en==1'b1)
			r_17_55 <= data_in;
	if (addr_selector[17]&addr_selector[56])
		data_out <= r_17_56;
		if (write_en==1'b1)
			r_17_56 <= data_in;
	if (addr_selector[17]&addr_selector[57])
		data_out <= r_17_57;
		if (write_en==1'b1)
			r_17_57 <= data_in;
	if (addr_selector[17]&addr_selector[58])
		data_out <= r_17_58;
		if (write_en==1'b1)
			r_17_58 <= data_in;
	if (addr_selector[17]&addr_selector[59])
		data_out <= r_17_59;
		if (write_en==1'b1)
			r_17_59 <= data_in;
	if (addr_selector[17]&addr_selector[60])
		data_out <= r_17_60;
		if (write_en==1'b1)
			r_17_60 <= data_in;
	if (addr_selector[17]&addr_selector[61])
		data_out <= r_17_61;
		if (write_en==1'b1)
			r_17_61 <= data_in;
	if (addr_selector[17]&addr_selector[62])
		data_out <= r_17_62;
		if (write_en==1'b1)
			r_17_62 <= data_in;
	if (addr_selector[17]&addr_selector[63])
		data_out <= r_17_63;
		if (write_en==1'b1)
			r_17_63 <= data_in;
	if (addr_selector[18]&addr_selector[0])
		data_out <= r_18_0;
		if (write_en==1'b1)
			r_18_0 <= data_in;
	if (addr_selector[18]&addr_selector[1])
		data_out <= r_18_1;
		if (write_en==1'b1)
			r_18_1 <= data_in;
	if (addr_selector[18]&addr_selector[2])
		data_out <= r_18_2;
		if (write_en==1'b1)
			r_18_2 <= data_in;
	if (addr_selector[18]&addr_selector[3])
		data_out <= r_18_3;
		if (write_en==1'b1)
			r_18_3 <= data_in;
	if (addr_selector[18]&addr_selector[4])
		data_out <= r_18_4;
		if (write_en==1'b1)
			r_18_4 <= data_in;
	if (addr_selector[18]&addr_selector[5])
		data_out <= r_18_5;
		if (write_en==1'b1)
			r_18_5 <= data_in;
	if (addr_selector[18]&addr_selector[6])
		data_out <= r_18_6;
		if (write_en==1'b1)
			r_18_6 <= data_in;
	if (addr_selector[18]&addr_selector[7])
		data_out <= r_18_7;
		if (write_en==1'b1)
			r_18_7 <= data_in;
	if (addr_selector[18]&addr_selector[8])
		data_out <= r_18_8;
		if (write_en==1'b1)
			r_18_8 <= data_in;
	if (addr_selector[18]&addr_selector[9])
		data_out <= r_18_9;
		if (write_en==1'b1)
			r_18_9 <= data_in;
	if (addr_selector[18]&addr_selector[10])
		data_out <= r_18_10;
		if (write_en==1'b1)
			r_18_10 <= data_in;
	if (addr_selector[18]&addr_selector[11])
		data_out <= r_18_11;
		if (write_en==1'b1)
			r_18_11 <= data_in;
	if (addr_selector[18]&addr_selector[12])
		data_out <= r_18_12;
		if (write_en==1'b1)
			r_18_12 <= data_in;
	if (addr_selector[18]&addr_selector[13])
		data_out <= r_18_13;
		if (write_en==1'b1)
			r_18_13 <= data_in;
	if (addr_selector[18]&addr_selector[14])
		data_out <= r_18_14;
		if (write_en==1'b1)
			r_18_14 <= data_in;
	if (addr_selector[18]&addr_selector[15])
		data_out <= r_18_15;
		if (write_en==1'b1)
			r_18_15 <= data_in;
	if (addr_selector[18]&addr_selector[16])
		data_out <= r_18_16;
		if (write_en==1'b1)
			r_18_16 <= data_in;
	if (addr_selector[18]&addr_selector[17])
		data_out <= r_18_17;
		if (write_en==1'b1)
			r_18_17 <= data_in;
	if (addr_selector[18]&addr_selector[18])
		data_out <= r_18_18;
		if (write_en==1'b1)
			r_18_18 <= data_in;
	if (addr_selector[18]&addr_selector[19])
		data_out <= r_18_19;
		if (write_en==1'b1)
			r_18_19 <= data_in;
	if (addr_selector[18]&addr_selector[20])
		data_out <= r_18_20;
		if (write_en==1'b1)
			r_18_20 <= data_in;
	if (addr_selector[18]&addr_selector[21])
		data_out <= r_18_21;
		if (write_en==1'b1)
			r_18_21 <= data_in;
	if (addr_selector[18]&addr_selector[22])
		data_out <= r_18_22;
		if (write_en==1'b1)
			r_18_22 <= data_in;
	if (addr_selector[18]&addr_selector[23])
		data_out <= r_18_23;
		if (write_en==1'b1)
			r_18_23 <= data_in;
	if (addr_selector[18]&addr_selector[24])
		data_out <= r_18_24;
		if (write_en==1'b1)
			r_18_24 <= data_in;
	if (addr_selector[18]&addr_selector[25])
		data_out <= r_18_25;
		if (write_en==1'b1)
			r_18_25 <= data_in;
	if (addr_selector[18]&addr_selector[26])
		data_out <= r_18_26;
		if (write_en==1'b1)
			r_18_26 <= data_in;
	if (addr_selector[18]&addr_selector[27])
		data_out <= r_18_27;
		if (write_en==1'b1)
			r_18_27 <= data_in;
	if (addr_selector[18]&addr_selector[28])
		data_out <= r_18_28;
		if (write_en==1'b1)
			r_18_28 <= data_in;
	if (addr_selector[18]&addr_selector[29])
		data_out <= r_18_29;
		if (write_en==1'b1)
			r_18_29 <= data_in;
	if (addr_selector[18]&addr_selector[30])
		data_out <= r_18_30;
		if (write_en==1'b1)
			r_18_30 <= data_in;
	if (addr_selector[18]&addr_selector[31])
		data_out <= r_18_31;
		if (write_en==1'b1)
			r_18_31 <= data_in;
	if (addr_selector[18]&addr_selector[32])
		data_out <= r_18_32;
		if (write_en==1'b1)
			r_18_32 <= data_in;
	if (addr_selector[18]&addr_selector[33])
		data_out <= r_18_33;
		if (write_en==1'b1)
			r_18_33 <= data_in;
	if (addr_selector[18]&addr_selector[34])
		data_out <= r_18_34;
		if (write_en==1'b1)
			r_18_34 <= data_in;
	if (addr_selector[18]&addr_selector[35])
		data_out <= r_18_35;
		if (write_en==1'b1)
			r_18_35 <= data_in;
	if (addr_selector[18]&addr_selector[36])
		data_out <= r_18_36;
		if (write_en==1'b1)
			r_18_36 <= data_in;
	if (addr_selector[18]&addr_selector[37])
		data_out <= r_18_37;
		if (write_en==1'b1)
			r_18_37 <= data_in;
	if (addr_selector[18]&addr_selector[38])
		data_out <= r_18_38;
		if (write_en==1'b1)
			r_18_38 <= data_in;
	if (addr_selector[18]&addr_selector[39])
		data_out <= r_18_39;
		if (write_en==1'b1)
			r_18_39 <= data_in;
	if (addr_selector[18]&addr_selector[40])
		data_out <= r_18_40;
		if (write_en==1'b1)
			r_18_40 <= data_in;
	if (addr_selector[18]&addr_selector[41])
		data_out <= r_18_41;
		if (write_en==1'b1)
			r_18_41 <= data_in;
	if (addr_selector[18]&addr_selector[42])
		data_out <= r_18_42;
		if (write_en==1'b1)
			r_18_42 <= data_in;
	if (addr_selector[18]&addr_selector[43])
		data_out <= r_18_43;
		if (write_en==1'b1)
			r_18_43 <= data_in;
	if (addr_selector[18]&addr_selector[44])
		data_out <= r_18_44;
		if (write_en==1'b1)
			r_18_44 <= data_in;
	if (addr_selector[18]&addr_selector[45])
		data_out <= r_18_45;
		if (write_en==1'b1)
			r_18_45 <= data_in;
	if (addr_selector[18]&addr_selector[46])
		data_out <= r_18_46;
		if (write_en==1'b1)
			r_18_46 <= data_in;
	if (addr_selector[18]&addr_selector[47])
		data_out <= r_18_47;
		if (write_en==1'b1)
			r_18_47 <= data_in;
	if (addr_selector[18]&addr_selector[48])
		data_out <= r_18_48;
		if (write_en==1'b1)
			r_18_48 <= data_in;
	if (addr_selector[18]&addr_selector[49])
		data_out <= r_18_49;
		if (write_en==1'b1)
			r_18_49 <= data_in;
	if (addr_selector[18]&addr_selector[50])
		data_out <= r_18_50;
		if (write_en==1'b1)
			r_18_50 <= data_in;
	if (addr_selector[18]&addr_selector[51])
		data_out <= r_18_51;
		if (write_en==1'b1)
			r_18_51 <= data_in;
	if (addr_selector[18]&addr_selector[52])
		data_out <= r_18_52;
		if (write_en==1'b1)
			r_18_52 <= data_in;
	if (addr_selector[18]&addr_selector[53])
		data_out <= r_18_53;
		if (write_en==1'b1)
			r_18_53 <= data_in;
	if (addr_selector[18]&addr_selector[54])
		data_out <= r_18_54;
		if (write_en==1'b1)
			r_18_54 <= data_in;
	if (addr_selector[18]&addr_selector[55])
		data_out <= r_18_55;
		if (write_en==1'b1)
			r_18_55 <= data_in;
	if (addr_selector[18]&addr_selector[56])
		data_out <= r_18_56;
		if (write_en==1'b1)
			r_18_56 <= data_in;
	if (addr_selector[18]&addr_selector[57])
		data_out <= r_18_57;
		if (write_en==1'b1)
			r_18_57 <= data_in;
	if (addr_selector[18]&addr_selector[58])
		data_out <= r_18_58;
		if (write_en==1'b1)
			r_18_58 <= data_in;
	if (addr_selector[18]&addr_selector[59])
		data_out <= r_18_59;
		if (write_en==1'b1)
			r_18_59 <= data_in;
	if (addr_selector[18]&addr_selector[60])
		data_out <= r_18_60;
		if (write_en==1'b1)
			r_18_60 <= data_in;
	if (addr_selector[18]&addr_selector[61])
		data_out <= r_18_61;
		if (write_en==1'b1)
			r_18_61 <= data_in;
	if (addr_selector[18]&addr_selector[62])
		data_out <= r_18_62;
		if (write_en==1'b1)
			r_18_62 <= data_in;
	if (addr_selector[18]&addr_selector[63])
		data_out <= r_18_63;
		if (write_en==1'b1)
			r_18_63 <= data_in;
	if (addr_selector[19]&addr_selector[0])
		data_out <= r_19_0;
		if (write_en==1'b1)
			r_19_0 <= data_in;
	if (addr_selector[19]&addr_selector[1])
		data_out <= r_19_1;
		if (write_en==1'b1)
			r_19_1 <= data_in;
	if (addr_selector[19]&addr_selector[2])
		data_out <= r_19_2;
		if (write_en==1'b1)
			r_19_2 <= data_in;
	if (addr_selector[19]&addr_selector[3])
		data_out <= r_19_3;
		if (write_en==1'b1)
			r_19_3 <= data_in;
	if (addr_selector[19]&addr_selector[4])
		data_out <= r_19_4;
		if (write_en==1'b1)
			r_19_4 <= data_in;
	if (addr_selector[19]&addr_selector[5])
		data_out <= r_19_5;
		if (write_en==1'b1)
			r_19_5 <= data_in;
	if (addr_selector[19]&addr_selector[6])
		data_out <= r_19_6;
		if (write_en==1'b1)
			r_19_6 <= data_in;
	if (addr_selector[19]&addr_selector[7])
		data_out <= r_19_7;
		if (write_en==1'b1)
			r_19_7 <= data_in;
	if (addr_selector[19]&addr_selector[8])
		data_out <= r_19_8;
		if (write_en==1'b1)
			r_19_8 <= data_in;
	if (addr_selector[19]&addr_selector[9])
		data_out <= r_19_9;
		if (write_en==1'b1)
			r_19_9 <= data_in;
	if (addr_selector[19]&addr_selector[10])
		data_out <= r_19_10;
		if (write_en==1'b1)
			r_19_10 <= data_in;
	if (addr_selector[19]&addr_selector[11])
		data_out <= r_19_11;
		if (write_en==1'b1)
			r_19_11 <= data_in;
	if (addr_selector[19]&addr_selector[12])
		data_out <= r_19_12;
		if (write_en==1'b1)
			r_19_12 <= data_in;
	if (addr_selector[19]&addr_selector[13])
		data_out <= r_19_13;
		if (write_en==1'b1)
			r_19_13 <= data_in;
	if (addr_selector[19]&addr_selector[14])
		data_out <= r_19_14;
		if (write_en==1'b1)
			r_19_14 <= data_in;
	if (addr_selector[19]&addr_selector[15])
		data_out <= r_19_15;
		if (write_en==1'b1)
			r_19_15 <= data_in;
	if (addr_selector[19]&addr_selector[16])
		data_out <= r_19_16;
		if (write_en==1'b1)
			r_19_16 <= data_in;
	if (addr_selector[19]&addr_selector[17])
		data_out <= r_19_17;
		if (write_en==1'b1)
			r_19_17 <= data_in;
	if (addr_selector[19]&addr_selector[18])
		data_out <= r_19_18;
		if (write_en==1'b1)
			r_19_18 <= data_in;
	if (addr_selector[19]&addr_selector[19])
		data_out <= r_19_19;
		if (write_en==1'b1)
			r_19_19 <= data_in;
	if (addr_selector[19]&addr_selector[20])
		data_out <= r_19_20;
		if (write_en==1'b1)
			r_19_20 <= data_in;
	if (addr_selector[19]&addr_selector[21])
		data_out <= r_19_21;
		if (write_en==1'b1)
			r_19_21 <= data_in;
	if (addr_selector[19]&addr_selector[22])
		data_out <= r_19_22;
		if (write_en==1'b1)
			r_19_22 <= data_in;
	if (addr_selector[19]&addr_selector[23])
		data_out <= r_19_23;
		if (write_en==1'b1)
			r_19_23 <= data_in;
	if (addr_selector[19]&addr_selector[24])
		data_out <= r_19_24;
		if (write_en==1'b1)
			r_19_24 <= data_in;
	if (addr_selector[19]&addr_selector[25])
		data_out <= r_19_25;
		if (write_en==1'b1)
			r_19_25 <= data_in;
	if (addr_selector[19]&addr_selector[26])
		data_out <= r_19_26;
		if (write_en==1'b1)
			r_19_26 <= data_in;
	if (addr_selector[19]&addr_selector[27])
		data_out <= r_19_27;
		if (write_en==1'b1)
			r_19_27 <= data_in;
	if (addr_selector[19]&addr_selector[28])
		data_out <= r_19_28;
		if (write_en==1'b1)
			r_19_28 <= data_in;
	if (addr_selector[19]&addr_selector[29])
		data_out <= r_19_29;
		if (write_en==1'b1)
			r_19_29 <= data_in;
	if (addr_selector[19]&addr_selector[30])
		data_out <= r_19_30;
		if (write_en==1'b1)
			r_19_30 <= data_in;
	if (addr_selector[19]&addr_selector[31])
		data_out <= r_19_31;
		if (write_en==1'b1)
			r_19_31 <= data_in;
	if (addr_selector[19]&addr_selector[32])
		data_out <= r_19_32;
		if (write_en==1'b1)
			r_19_32 <= data_in;
	if (addr_selector[19]&addr_selector[33])
		data_out <= r_19_33;
		if (write_en==1'b1)
			r_19_33 <= data_in;
	if (addr_selector[19]&addr_selector[34])
		data_out <= r_19_34;
		if (write_en==1'b1)
			r_19_34 <= data_in;
	if (addr_selector[19]&addr_selector[35])
		data_out <= r_19_35;
		if (write_en==1'b1)
			r_19_35 <= data_in;
	if (addr_selector[19]&addr_selector[36])
		data_out <= r_19_36;
		if (write_en==1'b1)
			r_19_36 <= data_in;
	if (addr_selector[19]&addr_selector[37])
		data_out <= r_19_37;
		if (write_en==1'b1)
			r_19_37 <= data_in;
	if (addr_selector[19]&addr_selector[38])
		data_out <= r_19_38;
		if (write_en==1'b1)
			r_19_38 <= data_in;
	if (addr_selector[19]&addr_selector[39])
		data_out <= r_19_39;
		if (write_en==1'b1)
			r_19_39 <= data_in;
	if (addr_selector[19]&addr_selector[40])
		data_out <= r_19_40;
		if (write_en==1'b1)
			r_19_40 <= data_in;
	if (addr_selector[19]&addr_selector[41])
		data_out <= r_19_41;
		if (write_en==1'b1)
			r_19_41 <= data_in;
	if (addr_selector[19]&addr_selector[42])
		data_out <= r_19_42;
		if (write_en==1'b1)
			r_19_42 <= data_in;
	if (addr_selector[19]&addr_selector[43])
		data_out <= r_19_43;
		if (write_en==1'b1)
			r_19_43 <= data_in;
	if (addr_selector[19]&addr_selector[44])
		data_out <= r_19_44;
		if (write_en==1'b1)
			r_19_44 <= data_in;
	if (addr_selector[19]&addr_selector[45])
		data_out <= r_19_45;
		if (write_en==1'b1)
			r_19_45 <= data_in;
	if (addr_selector[19]&addr_selector[46])
		data_out <= r_19_46;
		if (write_en==1'b1)
			r_19_46 <= data_in;
	if (addr_selector[19]&addr_selector[47])
		data_out <= r_19_47;
		if (write_en==1'b1)
			r_19_47 <= data_in;
	if (addr_selector[19]&addr_selector[48])
		data_out <= r_19_48;
		if (write_en==1'b1)
			r_19_48 <= data_in;
	if (addr_selector[19]&addr_selector[49])
		data_out <= r_19_49;
		if (write_en==1'b1)
			r_19_49 <= data_in;
	if (addr_selector[19]&addr_selector[50])
		data_out <= r_19_50;
		if (write_en==1'b1)
			r_19_50 <= data_in;
	if (addr_selector[19]&addr_selector[51])
		data_out <= r_19_51;
		if (write_en==1'b1)
			r_19_51 <= data_in;
	if (addr_selector[19]&addr_selector[52])
		data_out <= r_19_52;
		if (write_en==1'b1)
			r_19_52 <= data_in;
	if (addr_selector[19]&addr_selector[53])
		data_out <= r_19_53;
		if (write_en==1'b1)
			r_19_53 <= data_in;
	if (addr_selector[19]&addr_selector[54])
		data_out <= r_19_54;
		if (write_en==1'b1)
			r_19_54 <= data_in;
	if (addr_selector[19]&addr_selector[55])
		data_out <= r_19_55;
		if (write_en==1'b1)
			r_19_55 <= data_in;
	if (addr_selector[19]&addr_selector[56])
		data_out <= r_19_56;
		if (write_en==1'b1)
			r_19_56 <= data_in;
	if (addr_selector[19]&addr_selector[57])
		data_out <= r_19_57;
		if (write_en==1'b1)
			r_19_57 <= data_in;
	if (addr_selector[19]&addr_selector[58])
		data_out <= r_19_58;
		if (write_en==1'b1)
			r_19_58 <= data_in;
	if (addr_selector[19]&addr_selector[59])
		data_out <= r_19_59;
		if (write_en==1'b1)
			r_19_59 <= data_in;
	if (addr_selector[19]&addr_selector[60])
		data_out <= r_19_60;
		if (write_en==1'b1)
			r_19_60 <= data_in;
	if (addr_selector[19]&addr_selector[61])
		data_out <= r_19_61;
		if (write_en==1'b1)
			r_19_61 <= data_in;
	if (addr_selector[19]&addr_selector[62])
		data_out <= r_19_62;
		if (write_en==1'b1)
			r_19_62 <= data_in;
	if (addr_selector[19]&addr_selector[63])
		data_out <= r_19_63;
		if (write_en==1'b1)
			r_19_63 <= data_in;
	if (addr_selector[20]&addr_selector[0])
		data_out <= r_20_0;
		if (write_en==1'b1)
			r_20_0 <= data_in;
	if (addr_selector[20]&addr_selector[1])
		data_out <= r_20_1;
		if (write_en==1'b1)
			r_20_1 <= data_in;
	if (addr_selector[20]&addr_selector[2])
		data_out <= r_20_2;
		if (write_en==1'b1)
			r_20_2 <= data_in;
	if (addr_selector[20]&addr_selector[3])
		data_out <= r_20_3;
		if (write_en==1'b1)
			r_20_3 <= data_in;
	if (addr_selector[20]&addr_selector[4])
		data_out <= r_20_4;
		if (write_en==1'b1)
			r_20_4 <= data_in;
	if (addr_selector[20]&addr_selector[5])
		data_out <= r_20_5;
		if (write_en==1'b1)
			r_20_5 <= data_in;
	if (addr_selector[20]&addr_selector[6])
		data_out <= r_20_6;
		if (write_en==1'b1)
			r_20_6 <= data_in;
	if (addr_selector[20]&addr_selector[7])
		data_out <= r_20_7;
		if (write_en==1'b1)
			r_20_7 <= data_in;
	if (addr_selector[20]&addr_selector[8])
		data_out <= r_20_8;
		if (write_en==1'b1)
			r_20_8 <= data_in;
	if (addr_selector[20]&addr_selector[9])
		data_out <= r_20_9;
		if (write_en==1'b1)
			r_20_9 <= data_in;
	if (addr_selector[20]&addr_selector[10])
		data_out <= r_20_10;
		if (write_en==1'b1)
			r_20_10 <= data_in;
	if (addr_selector[20]&addr_selector[11])
		data_out <= r_20_11;
		if (write_en==1'b1)
			r_20_11 <= data_in;
	if (addr_selector[20]&addr_selector[12])
		data_out <= r_20_12;
		if (write_en==1'b1)
			r_20_12 <= data_in;
	if (addr_selector[20]&addr_selector[13])
		data_out <= r_20_13;
		if (write_en==1'b1)
			r_20_13 <= data_in;
	if (addr_selector[20]&addr_selector[14])
		data_out <= r_20_14;
		if (write_en==1'b1)
			r_20_14 <= data_in;
	if (addr_selector[20]&addr_selector[15])
		data_out <= r_20_15;
		if (write_en==1'b1)
			r_20_15 <= data_in;
	if (addr_selector[20]&addr_selector[16])
		data_out <= r_20_16;
		if (write_en==1'b1)
			r_20_16 <= data_in;
	if (addr_selector[20]&addr_selector[17])
		data_out <= r_20_17;
		if (write_en==1'b1)
			r_20_17 <= data_in;
	if (addr_selector[20]&addr_selector[18])
		data_out <= r_20_18;
		if (write_en==1'b1)
			r_20_18 <= data_in;
	if (addr_selector[20]&addr_selector[19])
		data_out <= r_20_19;
		if (write_en==1'b1)
			r_20_19 <= data_in;
	if (addr_selector[20]&addr_selector[20])
		data_out <= r_20_20;
		if (write_en==1'b1)
			r_20_20 <= data_in;
	if (addr_selector[20]&addr_selector[21])
		data_out <= r_20_21;
		if (write_en==1'b1)
			r_20_21 <= data_in;
	if (addr_selector[20]&addr_selector[22])
		data_out <= r_20_22;
		if (write_en==1'b1)
			r_20_22 <= data_in;
	if (addr_selector[20]&addr_selector[23])
		data_out <= r_20_23;
		if (write_en==1'b1)
			r_20_23 <= data_in;
	if (addr_selector[20]&addr_selector[24])
		data_out <= r_20_24;
		if (write_en==1'b1)
			r_20_24 <= data_in;
	if (addr_selector[20]&addr_selector[25])
		data_out <= r_20_25;
		if (write_en==1'b1)
			r_20_25 <= data_in;
	if (addr_selector[20]&addr_selector[26])
		data_out <= r_20_26;
		if (write_en==1'b1)
			r_20_26 <= data_in;
	if (addr_selector[20]&addr_selector[27])
		data_out <= r_20_27;
		if (write_en==1'b1)
			r_20_27 <= data_in;
	if (addr_selector[20]&addr_selector[28])
		data_out <= r_20_28;
		if (write_en==1'b1)
			r_20_28 <= data_in;
	if (addr_selector[20]&addr_selector[29])
		data_out <= r_20_29;
		if (write_en==1'b1)
			r_20_29 <= data_in;
	if (addr_selector[20]&addr_selector[30])
		data_out <= r_20_30;
		if (write_en==1'b1)
			r_20_30 <= data_in;
	if (addr_selector[20]&addr_selector[31])
		data_out <= r_20_31;
		if (write_en==1'b1)
			r_20_31 <= data_in;
	if (addr_selector[20]&addr_selector[32])
		data_out <= r_20_32;
		if (write_en==1'b1)
			r_20_32 <= data_in;
	if (addr_selector[20]&addr_selector[33])
		data_out <= r_20_33;
		if (write_en==1'b1)
			r_20_33 <= data_in;
	if (addr_selector[20]&addr_selector[34])
		data_out <= r_20_34;
		if (write_en==1'b1)
			r_20_34 <= data_in;
	if (addr_selector[20]&addr_selector[35])
		data_out <= r_20_35;
		if (write_en==1'b1)
			r_20_35 <= data_in;
	if (addr_selector[20]&addr_selector[36])
		data_out <= r_20_36;
		if (write_en==1'b1)
			r_20_36 <= data_in;
	if (addr_selector[20]&addr_selector[37])
		data_out <= r_20_37;
		if (write_en==1'b1)
			r_20_37 <= data_in;
	if (addr_selector[20]&addr_selector[38])
		data_out <= r_20_38;
		if (write_en==1'b1)
			r_20_38 <= data_in;
	if (addr_selector[20]&addr_selector[39])
		data_out <= r_20_39;
		if (write_en==1'b1)
			r_20_39 <= data_in;
	if (addr_selector[20]&addr_selector[40])
		data_out <= r_20_40;
		if (write_en==1'b1)
			r_20_40 <= data_in;
	if (addr_selector[20]&addr_selector[41])
		data_out <= r_20_41;
		if (write_en==1'b1)
			r_20_41 <= data_in;
	if (addr_selector[20]&addr_selector[42])
		data_out <= r_20_42;
		if (write_en==1'b1)
			r_20_42 <= data_in;
	if (addr_selector[20]&addr_selector[43])
		data_out <= r_20_43;
		if (write_en==1'b1)
			r_20_43 <= data_in;
	if (addr_selector[20]&addr_selector[44])
		data_out <= r_20_44;
		if (write_en==1'b1)
			r_20_44 <= data_in;
	if (addr_selector[20]&addr_selector[45])
		data_out <= r_20_45;
		if (write_en==1'b1)
			r_20_45 <= data_in;
	if (addr_selector[20]&addr_selector[46])
		data_out <= r_20_46;
		if (write_en==1'b1)
			r_20_46 <= data_in;
	if (addr_selector[20]&addr_selector[47])
		data_out <= r_20_47;
		if (write_en==1'b1)
			r_20_47 <= data_in;
	if (addr_selector[20]&addr_selector[48])
		data_out <= r_20_48;
		if (write_en==1'b1)
			r_20_48 <= data_in;
	if (addr_selector[20]&addr_selector[49])
		data_out <= r_20_49;
		if (write_en==1'b1)
			r_20_49 <= data_in;
	if (addr_selector[20]&addr_selector[50])
		data_out <= r_20_50;
		if (write_en==1'b1)
			r_20_50 <= data_in;
	if (addr_selector[20]&addr_selector[51])
		data_out <= r_20_51;
		if (write_en==1'b1)
			r_20_51 <= data_in;
	if (addr_selector[20]&addr_selector[52])
		data_out <= r_20_52;
		if (write_en==1'b1)
			r_20_52 <= data_in;
	if (addr_selector[20]&addr_selector[53])
		data_out <= r_20_53;
		if (write_en==1'b1)
			r_20_53 <= data_in;
	if (addr_selector[20]&addr_selector[54])
		data_out <= r_20_54;
		if (write_en==1'b1)
			r_20_54 <= data_in;
	if (addr_selector[20]&addr_selector[55])
		data_out <= r_20_55;
		if (write_en==1'b1)
			r_20_55 <= data_in;
	if (addr_selector[20]&addr_selector[56])
		data_out <= r_20_56;
		if (write_en==1'b1)
			r_20_56 <= data_in;
	if (addr_selector[20]&addr_selector[57])
		data_out <= r_20_57;
		if (write_en==1'b1)
			r_20_57 <= data_in;
	if (addr_selector[20]&addr_selector[58])
		data_out <= r_20_58;
		if (write_en==1'b1)
			r_20_58 <= data_in;
	if (addr_selector[20]&addr_selector[59])
		data_out <= r_20_59;
		if (write_en==1'b1)
			r_20_59 <= data_in;
	if (addr_selector[20]&addr_selector[60])
		data_out <= r_20_60;
		if (write_en==1'b1)
			r_20_60 <= data_in;
	if (addr_selector[20]&addr_selector[61])
		data_out <= r_20_61;
		if (write_en==1'b1)
			r_20_61 <= data_in;
	if (addr_selector[20]&addr_selector[62])
		data_out <= r_20_62;
		if (write_en==1'b1)
			r_20_62 <= data_in;
	if (addr_selector[20]&addr_selector[63])
		data_out <= r_20_63;
		if (write_en==1'b1)
			r_20_63 <= data_in;
	if (addr_selector[21]&addr_selector[0])
		data_out <= r_21_0;
		if (write_en==1'b1)
			r_21_0 <= data_in;
	if (addr_selector[21]&addr_selector[1])
		data_out <= r_21_1;
		if (write_en==1'b1)
			r_21_1 <= data_in;
	if (addr_selector[21]&addr_selector[2])
		data_out <= r_21_2;
		if (write_en==1'b1)
			r_21_2 <= data_in;
	if (addr_selector[21]&addr_selector[3])
		data_out <= r_21_3;
		if (write_en==1'b1)
			r_21_3 <= data_in;
	if (addr_selector[21]&addr_selector[4])
		data_out <= r_21_4;
		if (write_en==1'b1)
			r_21_4 <= data_in;
	if (addr_selector[21]&addr_selector[5])
		data_out <= r_21_5;
		if (write_en==1'b1)
			r_21_5 <= data_in;
	if (addr_selector[21]&addr_selector[6])
		data_out <= r_21_6;
		if (write_en==1'b1)
			r_21_6 <= data_in;
	if (addr_selector[21]&addr_selector[7])
		data_out <= r_21_7;
		if (write_en==1'b1)
			r_21_7 <= data_in;
	if (addr_selector[21]&addr_selector[8])
		data_out <= r_21_8;
		if (write_en==1'b1)
			r_21_8 <= data_in;
	if (addr_selector[21]&addr_selector[9])
		data_out <= r_21_9;
		if (write_en==1'b1)
			r_21_9 <= data_in;
	if (addr_selector[21]&addr_selector[10])
		data_out <= r_21_10;
		if (write_en==1'b1)
			r_21_10 <= data_in;
	if (addr_selector[21]&addr_selector[11])
		data_out <= r_21_11;
		if (write_en==1'b1)
			r_21_11 <= data_in;
	if (addr_selector[21]&addr_selector[12])
		data_out <= r_21_12;
		if (write_en==1'b1)
			r_21_12 <= data_in;
	if (addr_selector[21]&addr_selector[13])
		data_out <= r_21_13;
		if (write_en==1'b1)
			r_21_13 <= data_in;
	if (addr_selector[21]&addr_selector[14])
		data_out <= r_21_14;
		if (write_en==1'b1)
			r_21_14 <= data_in;
	if (addr_selector[21]&addr_selector[15])
		data_out <= r_21_15;
		if (write_en==1'b1)
			r_21_15 <= data_in;
	if (addr_selector[21]&addr_selector[16])
		data_out <= r_21_16;
		if (write_en==1'b1)
			r_21_16 <= data_in;
	if (addr_selector[21]&addr_selector[17])
		data_out <= r_21_17;
		if (write_en==1'b1)
			r_21_17 <= data_in;
	if (addr_selector[21]&addr_selector[18])
		data_out <= r_21_18;
		if (write_en==1'b1)
			r_21_18 <= data_in;
	if (addr_selector[21]&addr_selector[19])
		data_out <= r_21_19;
		if (write_en==1'b1)
			r_21_19 <= data_in;
	if (addr_selector[21]&addr_selector[20])
		data_out <= r_21_20;
		if (write_en==1'b1)
			r_21_20 <= data_in;
	if (addr_selector[21]&addr_selector[21])
		data_out <= r_21_21;
		if (write_en==1'b1)
			r_21_21 <= data_in;
	if (addr_selector[21]&addr_selector[22])
		data_out <= r_21_22;
		if (write_en==1'b1)
			r_21_22 <= data_in;
	if (addr_selector[21]&addr_selector[23])
		data_out <= r_21_23;
		if (write_en==1'b1)
			r_21_23 <= data_in;
	if (addr_selector[21]&addr_selector[24])
		data_out <= r_21_24;
		if (write_en==1'b1)
			r_21_24 <= data_in;
	if (addr_selector[21]&addr_selector[25])
		data_out <= r_21_25;
		if (write_en==1'b1)
			r_21_25 <= data_in;
	if (addr_selector[21]&addr_selector[26])
		data_out <= r_21_26;
		if (write_en==1'b1)
			r_21_26 <= data_in;
	if (addr_selector[21]&addr_selector[27])
		data_out <= r_21_27;
		if (write_en==1'b1)
			r_21_27 <= data_in;
	if (addr_selector[21]&addr_selector[28])
		data_out <= r_21_28;
		if (write_en==1'b1)
			r_21_28 <= data_in;
	if (addr_selector[21]&addr_selector[29])
		data_out <= r_21_29;
		if (write_en==1'b1)
			r_21_29 <= data_in;
	if (addr_selector[21]&addr_selector[30])
		data_out <= r_21_30;
		if (write_en==1'b1)
			r_21_30 <= data_in;
	if (addr_selector[21]&addr_selector[31])
		data_out <= r_21_31;
		if (write_en==1'b1)
			r_21_31 <= data_in;
	if (addr_selector[21]&addr_selector[32])
		data_out <= r_21_32;
		if (write_en==1'b1)
			r_21_32 <= data_in;
	if (addr_selector[21]&addr_selector[33])
		data_out <= r_21_33;
		if (write_en==1'b1)
			r_21_33 <= data_in;
	if (addr_selector[21]&addr_selector[34])
		data_out <= r_21_34;
		if (write_en==1'b1)
			r_21_34 <= data_in;
	if (addr_selector[21]&addr_selector[35])
		data_out <= r_21_35;
		if (write_en==1'b1)
			r_21_35 <= data_in;
	if (addr_selector[21]&addr_selector[36])
		data_out <= r_21_36;
		if (write_en==1'b1)
			r_21_36 <= data_in;
	if (addr_selector[21]&addr_selector[37])
		data_out <= r_21_37;
		if (write_en==1'b1)
			r_21_37 <= data_in;
	if (addr_selector[21]&addr_selector[38])
		data_out <= r_21_38;
		if (write_en==1'b1)
			r_21_38 <= data_in;
	if (addr_selector[21]&addr_selector[39])
		data_out <= r_21_39;
		if (write_en==1'b1)
			r_21_39 <= data_in;
	if (addr_selector[21]&addr_selector[40])
		data_out <= r_21_40;
		if (write_en==1'b1)
			r_21_40 <= data_in;
	if (addr_selector[21]&addr_selector[41])
		data_out <= r_21_41;
		if (write_en==1'b1)
			r_21_41 <= data_in;
	if (addr_selector[21]&addr_selector[42])
		data_out <= r_21_42;
		if (write_en==1'b1)
			r_21_42 <= data_in;
	if (addr_selector[21]&addr_selector[43])
		data_out <= r_21_43;
		if (write_en==1'b1)
			r_21_43 <= data_in;
	if (addr_selector[21]&addr_selector[44])
		data_out <= r_21_44;
		if (write_en==1'b1)
			r_21_44 <= data_in;
	if (addr_selector[21]&addr_selector[45])
		data_out <= r_21_45;
		if (write_en==1'b1)
			r_21_45 <= data_in;
	if (addr_selector[21]&addr_selector[46])
		data_out <= r_21_46;
		if (write_en==1'b1)
			r_21_46 <= data_in;
	if (addr_selector[21]&addr_selector[47])
		data_out <= r_21_47;
		if (write_en==1'b1)
			r_21_47 <= data_in;
	if (addr_selector[21]&addr_selector[48])
		data_out <= r_21_48;
		if (write_en==1'b1)
			r_21_48 <= data_in;
	if (addr_selector[21]&addr_selector[49])
		data_out <= r_21_49;
		if (write_en==1'b1)
			r_21_49 <= data_in;
	if (addr_selector[21]&addr_selector[50])
		data_out <= r_21_50;
		if (write_en==1'b1)
			r_21_50 <= data_in;
	if (addr_selector[21]&addr_selector[51])
		data_out <= r_21_51;
		if (write_en==1'b1)
			r_21_51 <= data_in;
	if (addr_selector[21]&addr_selector[52])
		data_out <= r_21_52;
		if (write_en==1'b1)
			r_21_52 <= data_in;
	if (addr_selector[21]&addr_selector[53])
		data_out <= r_21_53;
		if (write_en==1'b1)
			r_21_53 <= data_in;
	if (addr_selector[21]&addr_selector[54])
		data_out <= r_21_54;
		if (write_en==1'b1)
			r_21_54 <= data_in;
	if (addr_selector[21]&addr_selector[55])
		data_out <= r_21_55;
		if (write_en==1'b1)
			r_21_55 <= data_in;
	if (addr_selector[21]&addr_selector[56])
		data_out <= r_21_56;
		if (write_en==1'b1)
			r_21_56 <= data_in;
	if (addr_selector[21]&addr_selector[57])
		data_out <= r_21_57;
		if (write_en==1'b1)
			r_21_57 <= data_in;
	if (addr_selector[21]&addr_selector[58])
		data_out <= r_21_58;
		if (write_en==1'b1)
			r_21_58 <= data_in;
	if (addr_selector[21]&addr_selector[59])
		data_out <= r_21_59;
		if (write_en==1'b1)
			r_21_59 <= data_in;
	if (addr_selector[21]&addr_selector[60])
		data_out <= r_21_60;
		if (write_en==1'b1)
			r_21_60 <= data_in;
	if (addr_selector[21]&addr_selector[61])
		data_out <= r_21_61;
		if (write_en==1'b1)
			r_21_61 <= data_in;
	if (addr_selector[21]&addr_selector[62])
		data_out <= r_21_62;
		if (write_en==1'b1)
			r_21_62 <= data_in;
	if (addr_selector[21]&addr_selector[63])
		data_out <= r_21_63;
		if (write_en==1'b1)
			r_21_63 <= data_in;
	if (addr_selector[22]&addr_selector[0])
		data_out <= r_22_0;
		if (write_en==1'b1)
			r_22_0 <= data_in;
	if (addr_selector[22]&addr_selector[1])
		data_out <= r_22_1;
		if (write_en==1'b1)
			r_22_1 <= data_in;
	if (addr_selector[22]&addr_selector[2])
		data_out <= r_22_2;
		if (write_en==1'b1)
			r_22_2 <= data_in;
	if (addr_selector[22]&addr_selector[3])
		data_out <= r_22_3;
		if (write_en==1'b1)
			r_22_3 <= data_in;
	if (addr_selector[22]&addr_selector[4])
		data_out <= r_22_4;
		if (write_en==1'b1)
			r_22_4 <= data_in;
	if (addr_selector[22]&addr_selector[5])
		data_out <= r_22_5;
		if (write_en==1'b1)
			r_22_5 <= data_in;
	if (addr_selector[22]&addr_selector[6])
		data_out <= r_22_6;
		if (write_en==1'b1)
			r_22_6 <= data_in;
	if (addr_selector[22]&addr_selector[7])
		data_out <= r_22_7;
		if (write_en==1'b1)
			r_22_7 <= data_in;
	if (addr_selector[22]&addr_selector[8])
		data_out <= r_22_8;
		if (write_en==1'b1)
			r_22_8 <= data_in;
	if (addr_selector[22]&addr_selector[9])
		data_out <= r_22_9;
		if (write_en==1'b1)
			r_22_9 <= data_in;
	if (addr_selector[22]&addr_selector[10])
		data_out <= r_22_10;
		if (write_en==1'b1)
			r_22_10 <= data_in;
	if (addr_selector[22]&addr_selector[11])
		data_out <= r_22_11;
		if (write_en==1'b1)
			r_22_11 <= data_in;
	if (addr_selector[22]&addr_selector[12])
		data_out <= r_22_12;
		if (write_en==1'b1)
			r_22_12 <= data_in;
	if (addr_selector[22]&addr_selector[13])
		data_out <= r_22_13;
		if (write_en==1'b1)
			r_22_13 <= data_in;
	if (addr_selector[22]&addr_selector[14])
		data_out <= r_22_14;
		if (write_en==1'b1)
			r_22_14 <= data_in;
	if (addr_selector[22]&addr_selector[15])
		data_out <= r_22_15;
		if (write_en==1'b1)
			r_22_15 <= data_in;
	if (addr_selector[22]&addr_selector[16])
		data_out <= r_22_16;
		if (write_en==1'b1)
			r_22_16 <= data_in;
	if (addr_selector[22]&addr_selector[17])
		data_out <= r_22_17;
		if (write_en==1'b1)
			r_22_17 <= data_in;
	if (addr_selector[22]&addr_selector[18])
		data_out <= r_22_18;
		if (write_en==1'b1)
			r_22_18 <= data_in;
	if (addr_selector[22]&addr_selector[19])
		data_out <= r_22_19;
		if (write_en==1'b1)
			r_22_19 <= data_in;
	if (addr_selector[22]&addr_selector[20])
		data_out <= r_22_20;
		if (write_en==1'b1)
			r_22_20 <= data_in;
	if (addr_selector[22]&addr_selector[21])
		data_out <= r_22_21;
		if (write_en==1'b1)
			r_22_21 <= data_in;
	if (addr_selector[22]&addr_selector[22])
		data_out <= r_22_22;
		if (write_en==1'b1)
			r_22_22 <= data_in;
	if (addr_selector[22]&addr_selector[23])
		data_out <= r_22_23;
		if (write_en==1'b1)
			r_22_23 <= data_in;
	if (addr_selector[22]&addr_selector[24])
		data_out <= r_22_24;
		if (write_en==1'b1)
			r_22_24 <= data_in;
	if (addr_selector[22]&addr_selector[25])
		data_out <= r_22_25;
		if (write_en==1'b1)
			r_22_25 <= data_in;
	if (addr_selector[22]&addr_selector[26])
		data_out <= r_22_26;
		if (write_en==1'b1)
			r_22_26 <= data_in;
	if (addr_selector[22]&addr_selector[27])
		data_out <= r_22_27;
		if (write_en==1'b1)
			r_22_27 <= data_in;
	if (addr_selector[22]&addr_selector[28])
		data_out <= r_22_28;
		if (write_en==1'b1)
			r_22_28 <= data_in;
	if (addr_selector[22]&addr_selector[29])
		data_out <= r_22_29;
		if (write_en==1'b1)
			r_22_29 <= data_in;
	if (addr_selector[22]&addr_selector[30])
		data_out <= r_22_30;
		if (write_en==1'b1)
			r_22_30 <= data_in;
	if (addr_selector[22]&addr_selector[31])
		data_out <= r_22_31;
		if (write_en==1'b1)
			r_22_31 <= data_in;
	if (addr_selector[22]&addr_selector[32])
		data_out <= r_22_32;
		if (write_en==1'b1)
			r_22_32 <= data_in;
	if (addr_selector[22]&addr_selector[33])
		data_out <= r_22_33;
		if (write_en==1'b1)
			r_22_33 <= data_in;
	if (addr_selector[22]&addr_selector[34])
		data_out <= r_22_34;
		if (write_en==1'b1)
			r_22_34 <= data_in;
	if (addr_selector[22]&addr_selector[35])
		data_out <= r_22_35;
		if (write_en==1'b1)
			r_22_35 <= data_in;
	if (addr_selector[22]&addr_selector[36])
		data_out <= r_22_36;
		if (write_en==1'b1)
			r_22_36 <= data_in;
	if (addr_selector[22]&addr_selector[37])
		data_out <= r_22_37;
		if (write_en==1'b1)
			r_22_37 <= data_in;
	if (addr_selector[22]&addr_selector[38])
		data_out <= r_22_38;
		if (write_en==1'b1)
			r_22_38 <= data_in;
	if (addr_selector[22]&addr_selector[39])
		data_out <= r_22_39;
		if (write_en==1'b1)
			r_22_39 <= data_in;
	if (addr_selector[22]&addr_selector[40])
		data_out <= r_22_40;
		if (write_en==1'b1)
			r_22_40 <= data_in;
	if (addr_selector[22]&addr_selector[41])
		data_out <= r_22_41;
		if (write_en==1'b1)
			r_22_41 <= data_in;
	if (addr_selector[22]&addr_selector[42])
		data_out <= r_22_42;
		if (write_en==1'b1)
			r_22_42 <= data_in;
	if (addr_selector[22]&addr_selector[43])
		data_out <= r_22_43;
		if (write_en==1'b1)
			r_22_43 <= data_in;
	if (addr_selector[22]&addr_selector[44])
		data_out <= r_22_44;
		if (write_en==1'b1)
			r_22_44 <= data_in;
	if (addr_selector[22]&addr_selector[45])
		data_out <= r_22_45;
		if (write_en==1'b1)
			r_22_45 <= data_in;
	if (addr_selector[22]&addr_selector[46])
		data_out <= r_22_46;
		if (write_en==1'b1)
			r_22_46 <= data_in;
	if (addr_selector[22]&addr_selector[47])
		data_out <= r_22_47;
		if (write_en==1'b1)
			r_22_47 <= data_in;
	if (addr_selector[22]&addr_selector[48])
		data_out <= r_22_48;
		if (write_en==1'b1)
			r_22_48 <= data_in;
	if (addr_selector[22]&addr_selector[49])
		data_out <= r_22_49;
		if (write_en==1'b1)
			r_22_49 <= data_in;
	if (addr_selector[22]&addr_selector[50])
		data_out <= r_22_50;
		if (write_en==1'b1)
			r_22_50 <= data_in;
	if (addr_selector[22]&addr_selector[51])
		data_out <= r_22_51;
		if (write_en==1'b1)
			r_22_51 <= data_in;
	if (addr_selector[22]&addr_selector[52])
		data_out <= r_22_52;
		if (write_en==1'b1)
			r_22_52 <= data_in;
	if (addr_selector[22]&addr_selector[53])
		data_out <= r_22_53;
		if (write_en==1'b1)
			r_22_53 <= data_in;
	if (addr_selector[22]&addr_selector[54])
		data_out <= r_22_54;
		if (write_en==1'b1)
			r_22_54 <= data_in;
	if (addr_selector[22]&addr_selector[55])
		data_out <= r_22_55;
		if (write_en==1'b1)
			r_22_55 <= data_in;
	if (addr_selector[22]&addr_selector[56])
		data_out <= r_22_56;
		if (write_en==1'b1)
			r_22_56 <= data_in;
	if (addr_selector[22]&addr_selector[57])
		data_out <= r_22_57;
		if (write_en==1'b1)
			r_22_57 <= data_in;
	if (addr_selector[22]&addr_selector[58])
		data_out <= r_22_58;
		if (write_en==1'b1)
			r_22_58 <= data_in;
	if (addr_selector[22]&addr_selector[59])
		data_out <= r_22_59;
		if (write_en==1'b1)
			r_22_59 <= data_in;
	if (addr_selector[22]&addr_selector[60])
		data_out <= r_22_60;
		if (write_en==1'b1)
			r_22_60 <= data_in;
	if (addr_selector[22]&addr_selector[61])
		data_out <= r_22_61;
		if (write_en==1'b1)
			r_22_61 <= data_in;
	if (addr_selector[22]&addr_selector[62])
		data_out <= r_22_62;
		if (write_en==1'b1)
			r_22_62 <= data_in;
	if (addr_selector[22]&addr_selector[63])
		data_out <= r_22_63;
		if (write_en==1'b1)
			r_22_63 <= data_in;
	if (addr_selector[23]&addr_selector[0])
		data_out <= r_23_0;
		if (write_en==1'b1)
			r_23_0 <= data_in;
	if (addr_selector[23]&addr_selector[1])
		data_out <= r_23_1;
		if (write_en==1'b1)
			r_23_1 <= data_in;
	if (addr_selector[23]&addr_selector[2])
		data_out <= r_23_2;
		if (write_en==1'b1)
			r_23_2 <= data_in;
	if (addr_selector[23]&addr_selector[3])
		data_out <= r_23_3;
		if (write_en==1'b1)
			r_23_3 <= data_in;
	if (addr_selector[23]&addr_selector[4])
		data_out <= r_23_4;
		if (write_en==1'b1)
			r_23_4 <= data_in;
	if (addr_selector[23]&addr_selector[5])
		data_out <= r_23_5;
		if (write_en==1'b1)
			r_23_5 <= data_in;
	if (addr_selector[23]&addr_selector[6])
		data_out <= r_23_6;
		if (write_en==1'b1)
			r_23_6 <= data_in;
	if (addr_selector[23]&addr_selector[7])
		data_out <= r_23_7;
		if (write_en==1'b1)
			r_23_7 <= data_in;
	if (addr_selector[23]&addr_selector[8])
		data_out <= r_23_8;
		if (write_en==1'b1)
			r_23_8 <= data_in;
	if (addr_selector[23]&addr_selector[9])
		data_out <= r_23_9;
		if (write_en==1'b1)
			r_23_9 <= data_in;
	if (addr_selector[23]&addr_selector[10])
		data_out <= r_23_10;
		if (write_en==1'b1)
			r_23_10 <= data_in;
	if (addr_selector[23]&addr_selector[11])
		data_out <= r_23_11;
		if (write_en==1'b1)
			r_23_11 <= data_in;
	if (addr_selector[23]&addr_selector[12])
		data_out <= r_23_12;
		if (write_en==1'b1)
			r_23_12 <= data_in;
	if (addr_selector[23]&addr_selector[13])
		data_out <= r_23_13;
		if (write_en==1'b1)
			r_23_13 <= data_in;
	if (addr_selector[23]&addr_selector[14])
		data_out <= r_23_14;
		if (write_en==1'b1)
			r_23_14 <= data_in;
	if (addr_selector[23]&addr_selector[15])
		data_out <= r_23_15;
		if (write_en==1'b1)
			r_23_15 <= data_in;
	if (addr_selector[23]&addr_selector[16])
		data_out <= r_23_16;
		if (write_en==1'b1)
			r_23_16 <= data_in;
	if (addr_selector[23]&addr_selector[17])
		data_out <= r_23_17;
		if (write_en==1'b1)
			r_23_17 <= data_in;
	if (addr_selector[23]&addr_selector[18])
		data_out <= r_23_18;
		if (write_en==1'b1)
			r_23_18 <= data_in;
	if (addr_selector[23]&addr_selector[19])
		data_out <= r_23_19;
		if (write_en==1'b1)
			r_23_19 <= data_in;
	if (addr_selector[23]&addr_selector[20])
		data_out <= r_23_20;
		if (write_en==1'b1)
			r_23_20 <= data_in;
	if (addr_selector[23]&addr_selector[21])
		data_out <= r_23_21;
		if (write_en==1'b1)
			r_23_21 <= data_in;
	if (addr_selector[23]&addr_selector[22])
		data_out <= r_23_22;
		if (write_en==1'b1)
			r_23_22 <= data_in;
	if (addr_selector[23]&addr_selector[23])
		data_out <= r_23_23;
		if (write_en==1'b1)
			r_23_23 <= data_in;
	if (addr_selector[23]&addr_selector[24])
		data_out <= r_23_24;
		if (write_en==1'b1)
			r_23_24 <= data_in;
	if (addr_selector[23]&addr_selector[25])
		data_out <= r_23_25;
		if (write_en==1'b1)
			r_23_25 <= data_in;
	if (addr_selector[23]&addr_selector[26])
		data_out <= r_23_26;
		if (write_en==1'b1)
			r_23_26 <= data_in;
	if (addr_selector[23]&addr_selector[27])
		data_out <= r_23_27;
		if (write_en==1'b1)
			r_23_27 <= data_in;
	if (addr_selector[23]&addr_selector[28])
		data_out <= r_23_28;
		if (write_en==1'b1)
			r_23_28 <= data_in;
	if (addr_selector[23]&addr_selector[29])
		data_out <= r_23_29;
		if (write_en==1'b1)
			r_23_29 <= data_in;
	if (addr_selector[23]&addr_selector[30])
		data_out <= r_23_30;
		if (write_en==1'b1)
			r_23_30 <= data_in;
	if (addr_selector[23]&addr_selector[31])
		data_out <= r_23_31;
		if (write_en==1'b1)
			r_23_31 <= data_in;
	if (addr_selector[23]&addr_selector[32])
		data_out <= r_23_32;
		if (write_en==1'b1)
			r_23_32 <= data_in;
	if (addr_selector[23]&addr_selector[33])
		data_out <= r_23_33;
		if (write_en==1'b1)
			r_23_33 <= data_in;
	if (addr_selector[23]&addr_selector[34])
		data_out <= r_23_34;
		if (write_en==1'b1)
			r_23_34 <= data_in;
	if (addr_selector[23]&addr_selector[35])
		data_out <= r_23_35;
		if (write_en==1'b1)
			r_23_35 <= data_in;
	if (addr_selector[23]&addr_selector[36])
		data_out <= r_23_36;
		if (write_en==1'b1)
			r_23_36 <= data_in;
	if (addr_selector[23]&addr_selector[37])
		data_out <= r_23_37;
		if (write_en==1'b1)
			r_23_37 <= data_in;
	if (addr_selector[23]&addr_selector[38])
		data_out <= r_23_38;
		if (write_en==1'b1)
			r_23_38 <= data_in;
	if (addr_selector[23]&addr_selector[39])
		data_out <= r_23_39;
		if (write_en==1'b1)
			r_23_39 <= data_in;
	if (addr_selector[23]&addr_selector[40])
		data_out <= r_23_40;
		if (write_en==1'b1)
			r_23_40 <= data_in;
	if (addr_selector[23]&addr_selector[41])
		data_out <= r_23_41;
		if (write_en==1'b1)
			r_23_41 <= data_in;
	if (addr_selector[23]&addr_selector[42])
		data_out <= r_23_42;
		if (write_en==1'b1)
			r_23_42 <= data_in;
	if (addr_selector[23]&addr_selector[43])
		data_out <= r_23_43;
		if (write_en==1'b1)
			r_23_43 <= data_in;
	if (addr_selector[23]&addr_selector[44])
		data_out <= r_23_44;
		if (write_en==1'b1)
			r_23_44 <= data_in;
	if (addr_selector[23]&addr_selector[45])
		data_out <= r_23_45;
		if (write_en==1'b1)
			r_23_45 <= data_in;
	if (addr_selector[23]&addr_selector[46])
		data_out <= r_23_46;
		if (write_en==1'b1)
			r_23_46 <= data_in;
	if (addr_selector[23]&addr_selector[47])
		data_out <= r_23_47;
		if (write_en==1'b1)
			r_23_47 <= data_in;
	if (addr_selector[23]&addr_selector[48])
		data_out <= r_23_48;
		if (write_en==1'b1)
			r_23_48 <= data_in;
	if (addr_selector[23]&addr_selector[49])
		data_out <= r_23_49;
		if (write_en==1'b1)
			r_23_49 <= data_in;
	if (addr_selector[23]&addr_selector[50])
		data_out <= r_23_50;
		if (write_en==1'b1)
			r_23_50 <= data_in;
	if (addr_selector[23]&addr_selector[51])
		data_out <= r_23_51;
		if (write_en==1'b1)
			r_23_51 <= data_in;
	if (addr_selector[23]&addr_selector[52])
		data_out <= r_23_52;
		if (write_en==1'b1)
			r_23_52 <= data_in;
	if (addr_selector[23]&addr_selector[53])
		data_out <= r_23_53;
		if (write_en==1'b1)
			r_23_53 <= data_in;
	if (addr_selector[23]&addr_selector[54])
		data_out <= r_23_54;
		if (write_en==1'b1)
			r_23_54 <= data_in;
	if (addr_selector[23]&addr_selector[55])
		data_out <= r_23_55;
		if (write_en==1'b1)
			r_23_55 <= data_in;
	if (addr_selector[23]&addr_selector[56])
		data_out <= r_23_56;
		if (write_en==1'b1)
			r_23_56 <= data_in;
	if (addr_selector[23]&addr_selector[57])
		data_out <= r_23_57;
		if (write_en==1'b1)
			r_23_57 <= data_in;
	if (addr_selector[23]&addr_selector[58])
		data_out <= r_23_58;
		if (write_en==1'b1)
			r_23_58 <= data_in;
	if (addr_selector[23]&addr_selector[59])
		data_out <= r_23_59;
		if (write_en==1'b1)
			r_23_59 <= data_in;
	if (addr_selector[23]&addr_selector[60])
		data_out <= r_23_60;
		if (write_en==1'b1)
			r_23_60 <= data_in;
	if (addr_selector[23]&addr_selector[61])
		data_out <= r_23_61;
		if (write_en==1'b1)
			r_23_61 <= data_in;
	if (addr_selector[23]&addr_selector[62])
		data_out <= r_23_62;
		if (write_en==1'b1)
			r_23_62 <= data_in;
	if (addr_selector[23]&addr_selector[63])
		data_out <= r_23_63;
		if (write_en==1'b1)
			r_23_63 <= data_in;
	if (addr_selector[24]&addr_selector[0])
		data_out <= r_24_0;
		if (write_en==1'b1)
			r_24_0 <= data_in;
	if (addr_selector[24]&addr_selector[1])
		data_out <= r_24_1;
		if (write_en==1'b1)
			r_24_1 <= data_in;
	if (addr_selector[24]&addr_selector[2])
		data_out <= r_24_2;
		if (write_en==1'b1)
			r_24_2 <= data_in;
	if (addr_selector[24]&addr_selector[3])
		data_out <= r_24_3;
		if (write_en==1'b1)
			r_24_3 <= data_in;
	if (addr_selector[24]&addr_selector[4])
		data_out <= r_24_4;
		if (write_en==1'b1)
			r_24_4 <= data_in;
	if (addr_selector[24]&addr_selector[5])
		data_out <= r_24_5;
		if (write_en==1'b1)
			r_24_5 <= data_in;
	if (addr_selector[24]&addr_selector[6])
		data_out <= r_24_6;
		if (write_en==1'b1)
			r_24_6 <= data_in;
	if (addr_selector[24]&addr_selector[7])
		data_out <= r_24_7;
		if (write_en==1'b1)
			r_24_7 <= data_in;
	if (addr_selector[24]&addr_selector[8])
		data_out <= r_24_8;
		if (write_en==1'b1)
			r_24_8 <= data_in;
	if (addr_selector[24]&addr_selector[9])
		data_out <= r_24_9;
		if (write_en==1'b1)
			r_24_9 <= data_in;
	if (addr_selector[24]&addr_selector[10])
		data_out <= r_24_10;
		if (write_en==1'b1)
			r_24_10 <= data_in;
	if (addr_selector[24]&addr_selector[11])
		data_out <= r_24_11;
		if (write_en==1'b1)
			r_24_11 <= data_in;
	if (addr_selector[24]&addr_selector[12])
		data_out <= r_24_12;
		if (write_en==1'b1)
			r_24_12 <= data_in;
	if (addr_selector[24]&addr_selector[13])
		data_out <= r_24_13;
		if (write_en==1'b1)
			r_24_13 <= data_in;
	if (addr_selector[24]&addr_selector[14])
		data_out <= r_24_14;
		if (write_en==1'b1)
			r_24_14 <= data_in;
	if (addr_selector[24]&addr_selector[15])
		data_out <= r_24_15;
		if (write_en==1'b1)
			r_24_15 <= data_in;
	if (addr_selector[24]&addr_selector[16])
		data_out <= r_24_16;
		if (write_en==1'b1)
			r_24_16 <= data_in;
	if (addr_selector[24]&addr_selector[17])
		data_out <= r_24_17;
		if (write_en==1'b1)
			r_24_17 <= data_in;
	if (addr_selector[24]&addr_selector[18])
		data_out <= r_24_18;
		if (write_en==1'b1)
			r_24_18 <= data_in;
	if (addr_selector[24]&addr_selector[19])
		data_out <= r_24_19;
		if (write_en==1'b1)
			r_24_19 <= data_in;
	if (addr_selector[24]&addr_selector[20])
		data_out <= r_24_20;
		if (write_en==1'b1)
			r_24_20 <= data_in;
	if (addr_selector[24]&addr_selector[21])
		data_out <= r_24_21;
		if (write_en==1'b1)
			r_24_21 <= data_in;
	if (addr_selector[24]&addr_selector[22])
		data_out <= r_24_22;
		if (write_en==1'b1)
			r_24_22 <= data_in;
	if (addr_selector[24]&addr_selector[23])
		data_out <= r_24_23;
		if (write_en==1'b1)
			r_24_23 <= data_in;
	if (addr_selector[24]&addr_selector[24])
		data_out <= r_24_24;
		if (write_en==1'b1)
			r_24_24 <= data_in;
	if (addr_selector[24]&addr_selector[25])
		data_out <= r_24_25;
		if (write_en==1'b1)
			r_24_25 <= data_in;
	if (addr_selector[24]&addr_selector[26])
		data_out <= r_24_26;
		if (write_en==1'b1)
			r_24_26 <= data_in;
	if (addr_selector[24]&addr_selector[27])
		data_out <= r_24_27;
		if (write_en==1'b1)
			r_24_27 <= data_in;
	if (addr_selector[24]&addr_selector[28])
		data_out <= r_24_28;
		if (write_en==1'b1)
			r_24_28 <= data_in;
	if (addr_selector[24]&addr_selector[29])
		data_out <= r_24_29;
		if (write_en==1'b1)
			r_24_29 <= data_in;
	if (addr_selector[24]&addr_selector[30])
		data_out <= r_24_30;
		if (write_en==1'b1)
			r_24_30 <= data_in;
	if (addr_selector[24]&addr_selector[31])
		data_out <= r_24_31;
		if (write_en==1'b1)
			r_24_31 <= data_in;
	if (addr_selector[24]&addr_selector[32])
		data_out <= r_24_32;
		if (write_en==1'b1)
			r_24_32 <= data_in;
	if (addr_selector[24]&addr_selector[33])
		data_out <= r_24_33;
		if (write_en==1'b1)
			r_24_33 <= data_in;
	if (addr_selector[24]&addr_selector[34])
		data_out <= r_24_34;
		if (write_en==1'b1)
			r_24_34 <= data_in;
	if (addr_selector[24]&addr_selector[35])
		data_out <= r_24_35;
		if (write_en==1'b1)
			r_24_35 <= data_in;
	if (addr_selector[24]&addr_selector[36])
		data_out <= r_24_36;
		if (write_en==1'b1)
			r_24_36 <= data_in;
	if (addr_selector[24]&addr_selector[37])
		data_out <= r_24_37;
		if (write_en==1'b1)
			r_24_37 <= data_in;
	if (addr_selector[24]&addr_selector[38])
		data_out <= r_24_38;
		if (write_en==1'b1)
			r_24_38 <= data_in;
	if (addr_selector[24]&addr_selector[39])
		data_out <= r_24_39;
		if (write_en==1'b1)
			r_24_39 <= data_in;
	if (addr_selector[24]&addr_selector[40])
		data_out <= r_24_40;
		if (write_en==1'b1)
			r_24_40 <= data_in;
	if (addr_selector[24]&addr_selector[41])
		data_out <= r_24_41;
		if (write_en==1'b1)
			r_24_41 <= data_in;
	if (addr_selector[24]&addr_selector[42])
		data_out <= r_24_42;
		if (write_en==1'b1)
			r_24_42 <= data_in;
	if (addr_selector[24]&addr_selector[43])
		data_out <= r_24_43;
		if (write_en==1'b1)
			r_24_43 <= data_in;
	if (addr_selector[24]&addr_selector[44])
		data_out <= r_24_44;
		if (write_en==1'b1)
			r_24_44 <= data_in;
	if (addr_selector[24]&addr_selector[45])
		data_out <= r_24_45;
		if (write_en==1'b1)
			r_24_45 <= data_in;
	if (addr_selector[24]&addr_selector[46])
		data_out <= r_24_46;
		if (write_en==1'b1)
			r_24_46 <= data_in;
	if (addr_selector[24]&addr_selector[47])
		data_out <= r_24_47;
		if (write_en==1'b1)
			r_24_47 <= data_in;
	if (addr_selector[24]&addr_selector[48])
		data_out <= r_24_48;
		if (write_en==1'b1)
			r_24_48 <= data_in;
	if (addr_selector[24]&addr_selector[49])
		data_out <= r_24_49;
		if (write_en==1'b1)
			r_24_49 <= data_in;
	if (addr_selector[24]&addr_selector[50])
		data_out <= r_24_50;
		if (write_en==1'b1)
			r_24_50 <= data_in;
	if (addr_selector[24]&addr_selector[51])
		data_out <= r_24_51;
		if (write_en==1'b1)
			r_24_51 <= data_in;
	if (addr_selector[24]&addr_selector[52])
		data_out <= r_24_52;
		if (write_en==1'b1)
			r_24_52 <= data_in;
	if (addr_selector[24]&addr_selector[53])
		data_out <= r_24_53;
		if (write_en==1'b1)
			r_24_53 <= data_in;
	if (addr_selector[24]&addr_selector[54])
		data_out <= r_24_54;
		if (write_en==1'b1)
			r_24_54 <= data_in;
	if (addr_selector[24]&addr_selector[55])
		data_out <= r_24_55;
		if (write_en==1'b1)
			r_24_55 <= data_in;
	if (addr_selector[24]&addr_selector[56])
		data_out <= r_24_56;
		if (write_en==1'b1)
			r_24_56 <= data_in;
	if (addr_selector[24]&addr_selector[57])
		data_out <= r_24_57;
		if (write_en==1'b1)
			r_24_57 <= data_in;
	if (addr_selector[24]&addr_selector[58])
		data_out <= r_24_58;
		if (write_en==1'b1)
			r_24_58 <= data_in;
	if (addr_selector[24]&addr_selector[59])
		data_out <= r_24_59;
		if (write_en==1'b1)
			r_24_59 <= data_in;
	if (addr_selector[24]&addr_selector[60])
		data_out <= r_24_60;
		if (write_en==1'b1)
			r_24_60 <= data_in;
	if (addr_selector[24]&addr_selector[61])
		data_out <= r_24_61;
		if (write_en==1'b1)
			r_24_61 <= data_in;
	if (addr_selector[24]&addr_selector[62])
		data_out <= r_24_62;
		if (write_en==1'b1)
			r_24_62 <= data_in;
	if (addr_selector[24]&addr_selector[63])
		data_out <= r_24_63;
		if (write_en==1'b1)
			r_24_63 <= data_in;
	if (addr_selector[25]&addr_selector[0])
		data_out <= r_25_0;
		if (write_en==1'b1)
			r_25_0 <= data_in;
	if (addr_selector[25]&addr_selector[1])
		data_out <= r_25_1;
		if (write_en==1'b1)
			r_25_1 <= data_in;
	if (addr_selector[25]&addr_selector[2])
		data_out <= r_25_2;
		if (write_en==1'b1)
			r_25_2 <= data_in;
	if (addr_selector[25]&addr_selector[3])
		data_out <= r_25_3;
		if (write_en==1'b1)
			r_25_3 <= data_in;
	if (addr_selector[25]&addr_selector[4])
		data_out <= r_25_4;
		if (write_en==1'b1)
			r_25_4 <= data_in;
	if (addr_selector[25]&addr_selector[5])
		data_out <= r_25_5;
		if (write_en==1'b1)
			r_25_5 <= data_in;
	if (addr_selector[25]&addr_selector[6])
		data_out <= r_25_6;
		if (write_en==1'b1)
			r_25_6 <= data_in;
	if (addr_selector[25]&addr_selector[7])
		data_out <= r_25_7;
		if (write_en==1'b1)
			r_25_7 <= data_in;
	if (addr_selector[25]&addr_selector[8])
		data_out <= r_25_8;
		if (write_en==1'b1)
			r_25_8 <= data_in;
	if (addr_selector[25]&addr_selector[9])
		data_out <= r_25_9;
		if (write_en==1'b1)
			r_25_9 <= data_in;
	if (addr_selector[25]&addr_selector[10])
		data_out <= r_25_10;
		if (write_en==1'b1)
			r_25_10 <= data_in;
	if (addr_selector[25]&addr_selector[11])
		data_out <= r_25_11;
		if (write_en==1'b1)
			r_25_11 <= data_in;
	if (addr_selector[25]&addr_selector[12])
		data_out <= r_25_12;
		if (write_en==1'b1)
			r_25_12 <= data_in;
	if (addr_selector[25]&addr_selector[13])
		data_out <= r_25_13;
		if (write_en==1'b1)
			r_25_13 <= data_in;
	if (addr_selector[25]&addr_selector[14])
		data_out <= r_25_14;
		if (write_en==1'b1)
			r_25_14 <= data_in;
	if (addr_selector[25]&addr_selector[15])
		data_out <= r_25_15;
		if (write_en==1'b1)
			r_25_15 <= data_in;
	if (addr_selector[25]&addr_selector[16])
		data_out <= r_25_16;
		if (write_en==1'b1)
			r_25_16 <= data_in;
	if (addr_selector[25]&addr_selector[17])
		data_out <= r_25_17;
		if (write_en==1'b1)
			r_25_17 <= data_in;
	if (addr_selector[25]&addr_selector[18])
		data_out <= r_25_18;
		if (write_en==1'b1)
			r_25_18 <= data_in;
	if (addr_selector[25]&addr_selector[19])
		data_out <= r_25_19;
		if (write_en==1'b1)
			r_25_19 <= data_in;
	if (addr_selector[25]&addr_selector[20])
		data_out <= r_25_20;
		if (write_en==1'b1)
			r_25_20 <= data_in;
	if (addr_selector[25]&addr_selector[21])
		data_out <= r_25_21;
		if (write_en==1'b1)
			r_25_21 <= data_in;
	if (addr_selector[25]&addr_selector[22])
		data_out <= r_25_22;
		if (write_en==1'b1)
			r_25_22 <= data_in;
	if (addr_selector[25]&addr_selector[23])
		data_out <= r_25_23;
		if (write_en==1'b1)
			r_25_23 <= data_in;
	if (addr_selector[25]&addr_selector[24])
		data_out <= r_25_24;
		if (write_en==1'b1)
			r_25_24 <= data_in;
	if (addr_selector[25]&addr_selector[25])
		data_out <= r_25_25;
		if (write_en==1'b1)
			r_25_25 <= data_in;
	if (addr_selector[25]&addr_selector[26])
		data_out <= r_25_26;
		if (write_en==1'b1)
			r_25_26 <= data_in;
	if (addr_selector[25]&addr_selector[27])
		data_out <= r_25_27;
		if (write_en==1'b1)
			r_25_27 <= data_in;
	if (addr_selector[25]&addr_selector[28])
		data_out <= r_25_28;
		if (write_en==1'b1)
			r_25_28 <= data_in;
	if (addr_selector[25]&addr_selector[29])
		data_out <= r_25_29;
		if (write_en==1'b1)
			r_25_29 <= data_in;
	if (addr_selector[25]&addr_selector[30])
		data_out <= r_25_30;
		if (write_en==1'b1)
			r_25_30 <= data_in;
	if (addr_selector[25]&addr_selector[31])
		data_out <= r_25_31;
		if (write_en==1'b1)
			r_25_31 <= data_in;
	if (addr_selector[25]&addr_selector[32])
		data_out <= r_25_32;
		if (write_en==1'b1)
			r_25_32 <= data_in;
	if (addr_selector[25]&addr_selector[33])
		data_out <= r_25_33;
		if (write_en==1'b1)
			r_25_33 <= data_in;
	if (addr_selector[25]&addr_selector[34])
		data_out <= r_25_34;
		if (write_en==1'b1)
			r_25_34 <= data_in;
	if (addr_selector[25]&addr_selector[35])
		data_out <= r_25_35;
		if (write_en==1'b1)
			r_25_35 <= data_in;
	if (addr_selector[25]&addr_selector[36])
		data_out <= r_25_36;
		if (write_en==1'b1)
			r_25_36 <= data_in;
	if (addr_selector[25]&addr_selector[37])
		data_out <= r_25_37;
		if (write_en==1'b1)
			r_25_37 <= data_in;
	if (addr_selector[25]&addr_selector[38])
		data_out <= r_25_38;
		if (write_en==1'b1)
			r_25_38 <= data_in;
	if (addr_selector[25]&addr_selector[39])
		data_out <= r_25_39;
		if (write_en==1'b1)
			r_25_39 <= data_in;
	if (addr_selector[25]&addr_selector[40])
		data_out <= r_25_40;
		if (write_en==1'b1)
			r_25_40 <= data_in;
	if (addr_selector[25]&addr_selector[41])
		data_out <= r_25_41;
		if (write_en==1'b1)
			r_25_41 <= data_in;
	if (addr_selector[25]&addr_selector[42])
		data_out <= r_25_42;
		if (write_en==1'b1)
			r_25_42 <= data_in;
	if (addr_selector[25]&addr_selector[43])
		data_out <= r_25_43;
		if (write_en==1'b1)
			r_25_43 <= data_in;
	if (addr_selector[25]&addr_selector[44])
		data_out <= r_25_44;
		if (write_en==1'b1)
			r_25_44 <= data_in;
	if (addr_selector[25]&addr_selector[45])
		data_out <= r_25_45;
		if (write_en==1'b1)
			r_25_45 <= data_in;
	if (addr_selector[25]&addr_selector[46])
		data_out <= r_25_46;
		if (write_en==1'b1)
			r_25_46 <= data_in;
	if (addr_selector[25]&addr_selector[47])
		data_out <= r_25_47;
		if (write_en==1'b1)
			r_25_47 <= data_in;
	if (addr_selector[25]&addr_selector[48])
		data_out <= r_25_48;
		if (write_en==1'b1)
			r_25_48 <= data_in;
	if (addr_selector[25]&addr_selector[49])
		data_out <= r_25_49;
		if (write_en==1'b1)
			r_25_49 <= data_in;
	if (addr_selector[25]&addr_selector[50])
		data_out <= r_25_50;
		if (write_en==1'b1)
			r_25_50 <= data_in;
	if (addr_selector[25]&addr_selector[51])
		data_out <= r_25_51;
		if (write_en==1'b1)
			r_25_51 <= data_in;
	if (addr_selector[25]&addr_selector[52])
		data_out <= r_25_52;
		if (write_en==1'b1)
			r_25_52 <= data_in;
	if (addr_selector[25]&addr_selector[53])
		data_out <= r_25_53;
		if (write_en==1'b1)
			r_25_53 <= data_in;
	if (addr_selector[25]&addr_selector[54])
		data_out <= r_25_54;
		if (write_en==1'b1)
			r_25_54 <= data_in;
	if (addr_selector[25]&addr_selector[55])
		data_out <= r_25_55;
		if (write_en==1'b1)
			r_25_55 <= data_in;
	if (addr_selector[25]&addr_selector[56])
		data_out <= r_25_56;
		if (write_en==1'b1)
			r_25_56 <= data_in;
	if (addr_selector[25]&addr_selector[57])
		data_out <= r_25_57;
		if (write_en==1'b1)
			r_25_57 <= data_in;
	if (addr_selector[25]&addr_selector[58])
		data_out <= r_25_58;
		if (write_en==1'b1)
			r_25_58 <= data_in;
	if (addr_selector[25]&addr_selector[59])
		data_out <= r_25_59;
		if (write_en==1'b1)
			r_25_59 <= data_in;
	if (addr_selector[25]&addr_selector[60])
		data_out <= r_25_60;
		if (write_en==1'b1)
			r_25_60 <= data_in;
	if (addr_selector[25]&addr_selector[61])
		data_out <= r_25_61;
		if (write_en==1'b1)
			r_25_61 <= data_in;
	if (addr_selector[25]&addr_selector[62])
		data_out <= r_25_62;
		if (write_en==1'b1)
			r_25_62 <= data_in;
	if (addr_selector[25]&addr_selector[63])
		data_out <= r_25_63;
		if (write_en==1'b1)
			r_25_63 <= data_in;
	if (addr_selector[26]&addr_selector[0])
		data_out <= r_26_0;
		if (write_en==1'b1)
			r_26_0 <= data_in;
	if (addr_selector[26]&addr_selector[1])
		data_out <= r_26_1;
		if (write_en==1'b1)
			r_26_1 <= data_in;
	if (addr_selector[26]&addr_selector[2])
		data_out <= r_26_2;
		if (write_en==1'b1)
			r_26_2 <= data_in;
	if (addr_selector[26]&addr_selector[3])
		data_out <= r_26_3;
		if (write_en==1'b1)
			r_26_3 <= data_in;
	if (addr_selector[26]&addr_selector[4])
		data_out <= r_26_4;
		if (write_en==1'b1)
			r_26_4 <= data_in;
	if (addr_selector[26]&addr_selector[5])
		data_out <= r_26_5;
		if (write_en==1'b1)
			r_26_5 <= data_in;
	if (addr_selector[26]&addr_selector[6])
		data_out <= r_26_6;
		if (write_en==1'b1)
			r_26_6 <= data_in;
	if (addr_selector[26]&addr_selector[7])
		data_out <= r_26_7;
		if (write_en==1'b1)
			r_26_7 <= data_in;
	if (addr_selector[26]&addr_selector[8])
		data_out <= r_26_8;
		if (write_en==1'b1)
			r_26_8 <= data_in;
	if (addr_selector[26]&addr_selector[9])
		data_out <= r_26_9;
		if (write_en==1'b1)
			r_26_9 <= data_in;
	if (addr_selector[26]&addr_selector[10])
		data_out <= r_26_10;
		if (write_en==1'b1)
			r_26_10 <= data_in;
	if (addr_selector[26]&addr_selector[11])
		data_out <= r_26_11;
		if (write_en==1'b1)
			r_26_11 <= data_in;
	if (addr_selector[26]&addr_selector[12])
		data_out <= r_26_12;
		if (write_en==1'b1)
			r_26_12 <= data_in;
	if (addr_selector[26]&addr_selector[13])
		data_out <= r_26_13;
		if (write_en==1'b1)
			r_26_13 <= data_in;
	if (addr_selector[26]&addr_selector[14])
		data_out <= r_26_14;
		if (write_en==1'b1)
			r_26_14 <= data_in;
	if (addr_selector[26]&addr_selector[15])
		data_out <= r_26_15;
		if (write_en==1'b1)
			r_26_15 <= data_in;
	if (addr_selector[26]&addr_selector[16])
		data_out <= r_26_16;
		if (write_en==1'b1)
			r_26_16 <= data_in;
	if (addr_selector[26]&addr_selector[17])
		data_out <= r_26_17;
		if (write_en==1'b1)
			r_26_17 <= data_in;
	if (addr_selector[26]&addr_selector[18])
		data_out <= r_26_18;
		if (write_en==1'b1)
			r_26_18 <= data_in;
	if (addr_selector[26]&addr_selector[19])
		data_out <= r_26_19;
		if (write_en==1'b1)
			r_26_19 <= data_in;
	if (addr_selector[26]&addr_selector[20])
		data_out <= r_26_20;
		if (write_en==1'b1)
			r_26_20 <= data_in;
	if (addr_selector[26]&addr_selector[21])
		data_out <= r_26_21;
		if (write_en==1'b1)
			r_26_21 <= data_in;
	if (addr_selector[26]&addr_selector[22])
		data_out <= r_26_22;
		if (write_en==1'b1)
			r_26_22 <= data_in;
	if (addr_selector[26]&addr_selector[23])
		data_out <= r_26_23;
		if (write_en==1'b1)
			r_26_23 <= data_in;
	if (addr_selector[26]&addr_selector[24])
		data_out <= r_26_24;
		if (write_en==1'b1)
			r_26_24 <= data_in;
	if (addr_selector[26]&addr_selector[25])
		data_out <= r_26_25;
		if (write_en==1'b1)
			r_26_25 <= data_in;
	if (addr_selector[26]&addr_selector[26])
		data_out <= r_26_26;
		if (write_en==1'b1)
			r_26_26 <= data_in;
	if (addr_selector[26]&addr_selector[27])
		data_out <= r_26_27;
		if (write_en==1'b1)
			r_26_27 <= data_in;
	if (addr_selector[26]&addr_selector[28])
		data_out <= r_26_28;
		if (write_en==1'b1)
			r_26_28 <= data_in;
	if (addr_selector[26]&addr_selector[29])
		data_out <= r_26_29;
		if (write_en==1'b1)
			r_26_29 <= data_in;
	if (addr_selector[26]&addr_selector[30])
		data_out <= r_26_30;
		if (write_en==1'b1)
			r_26_30 <= data_in;
	if (addr_selector[26]&addr_selector[31])
		data_out <= r_26_31;
		if (write_en==1'b1)
			r_26_31 <= data_in;
	if (addr_selector[26]&addr_selector[32])
		data_out <= r_26_32;
		if (write_en==1'b1)
			r_26_32 <= data_in;
	if (addr_selector[26]&addr_selector[33])
		data_out <= r_26_33;
		if (write_en==1'b1)
			r_26_33 <= data_in;
	if (addr_selector[26]&addr_selector[34])
		data_out <= r_26_34;
		if (write_en==1'b1)
			r_26_34 <= data_in;
	if (addr_selector[26]&addr_selector[35])
		data_out <= r_26_35;
		if (write_en==1'b1)
			r_26_35 <= data_in;
	if (addr_selector[26]&addr_selector[36])
		data_out <= r_26_36;
		if (write_en==1'b1)
			r_26_36 <= data_in;
	if (addr_selector[26]&addr_selector[37])
		data_out <= r_26_37;
		if (write_en==1'b1)
			r_26_37 <= data_in;
	if (addr_selector[26]&addr_selector[38])
		data_out <= r_26_38;
		if (write_en==1'b1)
			r_26_38 <= data_in;
	if (addr_selector[26]&addr_selector[39])
		data_out <= r_26_39;
		if (write_en==1'b1)
			r_26_39 <= data_in;
	if (addr_selector[26]&addr_selector[40])
		data_out <= r_26_40;
		if (write_en==1'b1)
			r_26_40 <= data_in;
	if (addr_selector[26]&addr_selector[41])
		data_out <= r_26_41;
		if (write_en==1'b1)
			r_26_41 <= data_in;
	if (addr_selector[26]&addr_selector[42])
		data_out <= r_26_42;
		if (write_en==1'b1)
			r_26_42 <= data_in;
	if (addr_selector[26]&addr_selector[43])
		data_out <= r_26_43;
		if (write_en==1'b1)
			r_26_43 <= data_in;
	if (addr_selector[26]&addr_selector[44])
		data_out <= r_26_44;
		if (write_en==1'b1)
			r_26_44 <= data_in;
	if (addr_selector[26]&addr_selector[45])
		data_out <= r_26_45;
		if (write_en==1'b1)
			r_26_45 <= data_in;
	if (addr_selector[26]&addr_selector[46])
		data_out <= r_26_46;
		if (write_en==1'b1)
			r_26_46 <= data_in;
	if (addr_selector[26]&addr_selector[47])
		data_out <= r_26_47;
		if (write_en==1'b1)
			r_26_47 <= data_in;
	if (addr_selector[26]&addr_selector[48])
		data_out <= r_26_48;
		if (write_en==1'b1)
			r_26_48 <= data_in;
	if (addr_selector[26]&addr_selector[49])
		data_out <= r_26_49;
		if (write_en==1'b1)
			r_26_49 <= data_in;
	if (addr_selector[26]&addr_selector[50])
		data_out <= r_26_50;
		if (write_en==1'b1)
			r_26_50 <= data_in;
	if (addr_selector[26]&addr_selector[51])
		data_out <= r_26_51;
		if (write_en==1'b1)
			r_26_51 <= data_in;
	if (addr_selector[26]&addr_selector[52])
		data_out <= r_26_52;
		if (write_en==1'b1)
			r_26_52 <= data_in;
	if (addr_selector[26]&addr_selector[53])
		data_out <= r_26_53;
		if (write_en==1'b1)
			r_26_53 <= data_in;
	if (addr_selector[26]&addr_selector[54])
		data_out <= r_26_54;
		if (write_en==1'b1)
			r_26_54 <= data_in;
	if (addr_selector[26]&addr_selector[55])
		data_out <= r_26_55;
		if (write_en==1'b1)
			r_26_55 <= data_in;
	if (addr_selector[26]&addr_selector[56])
		data_out <= r_26_56;
		if (write_en==1'b1)
			r_26_56 <= data_in;
	if (addr_selector[26]&addr_selector[57])
		data_out <= r_26_57;
		if (write_en==1'b1)
			r_26_57 <= data_in;
	if (addr_selector[26]&addr_selector[58])
		data_out <= r_26_58;
		if (write_en==1'b1)
			r_26_58 <= data_in;
	if (addr_selector[26]&addr_selector[59])
		data_out <= r_26_59;
		if (write_en==1'b1)
			r_26_59 <= data_in;
	if (addr_selector[26]&addr_selector[60])
		data_out <= r_26_60;
		if (write_en==1'b1)
			r_26_60 <= data_in;
	if (addr_selector[26]&addr_selector[61])
		data_out <= r_26_61;
		if (write_en==1'b1)
			r_26_61 <= data_in;
	if (addr_selector[26]&addr_selector[62])
		data_out <= r_26_62;
		if (write_en==1'b1)
			r_26_62 <= data_in;
	if (addr_selector[26]&addr_selector[63])
		data_out <= r_26_63;
		if (write_en==1'b1)
			r_26_63 <= data_in;
	if (addr_selector[27]&addr_selector[0])
		data_out <= r_27_0;
		if (write_en==1'b1)
			r_27_0 <= data_in;
	if (addr_selector[27]&addr_selector[1])
		data_out <= r_27_1;
		if (write_en==1'b1)
			r_27_1 <= data_in;
	if (addr_selector[27]&addr_selector[2])
		data_out <= r_27_2;
		if (write_en==1'b1)
			r_27_2 <= data_in;
	if (addr_selector[27]&addr_selector[3])
		data_out <= r_27_3;
		if (write_en==1'b1)
			r_27_3 <= data_in;
	if (addr_selector[27]&addr_selector[4])
		data_out <= r_27_4;
		if (write_en==1'b1)
			r_27_4 <= data_in;
	if (addr_selector[27]&addr_selector[5])
		data_out <= r_27_5;
		if (write_en==1'b1)
			r_27_5 <= data_in;
	if (addr_selector[27]&addr_selector[6])
		data_out <= r_27_6;
		if (write_en==1'b1)
			r_27_6 <= data_in;
	if (addr_selector[27]&addr_selector[7])
		data_out <= r_27_7;
		if (write_en==1'b1)
			r_27_7 <= data_in;
	if (addr_selector[27]&addr_selector[8])
		data_out <= r_27_8;
		if (write_en==1'b1)
			r_27_8 <= data_in;
	if (addr_selector[27]&addr_selector[9])
		data_out <= r_27_9;
		if (write_en==1'b1)
			r_27_9 <= data_in;
	if (addr_selector[27]&addr_selector[10])
		data_out <= r_27_10;
		if (write_en==1'b1)
			r_27_10 <= data_in;
	if (addr_selector[27]&addr_selector[11])
		data_out <= r_27_11;
		if (write_en==1'b1)
			r_27_11 <= data_in;
	if (addr_selector[27]&addr_selector[12])
		data_out <= r_27_12;
		if (write_en==1'b1)
			r_27_12 <= data_in;
	if (addr_selector[27]&addr_selector[13])
		data_out <= r_27_13;
		if (write_en==1'b1)
			r_27_13 <= data_in;
	if (addr_selector[27]&addr_selector[14])
		data_out <= r_27_14;
		if (write_en==1'b1)
			r_27_14 <= data_in;
	if (addr_selector[27]&addr_selector[15])
		data_out <= r_27_15;
		if (write_en==1'b1)
			r_27_15 <= data_in;
	if (addr_selector[27]&addr_selector[16])
		data_out <= r_27_16;
		if (write_en==1'b1)
			r_27_16 <= data_in;
	if (addr_selector[27]&addr_selector[17])
		data_out <= r_27_17;
		if (write_en==1'b1)
			r_27_17 <= data_in;
	if (addr_selector[27]&addr_selector[18])
		data_out <= r_27_18;
		if (write_en==1'b1)
			r_27_18 <= data_in;
	if (addr_selector[27]&addr_selector[19])
		data_out <= r_27_19;
		if (write_en==1'b1)
			r_27_19 <= data_in;
	if (addr_selector[27]&addr_selector[20])
		data_out <= r_27_20;
		if (write_en==1'b1)
			r_27_20 <= data_in;
	if (addr_selector[27]&addr_selector[21])
		data_out <= r_27_21;
		if (write_en==1'b1)
			r_27_21 <= data_in;
	if (addr_selector[27]&addr_selector[22])
		data_out <= r_27_22;
		if (write_en==1'b1)
			r_27_22 <= data_in;
	if (addr_selector[27]&addr_selector[23])
		data_out <= r_27_23;
		if (write_en==1'b1)
			r_27_23 <= data_in;
	if (addr_selector[27]&addr_selector[24])
		data_out <= r_27_24;
		if (write_en==1'b1)
			r_27_24 <= data_in;
	if (addr_selector[27]&addr_selector[25])
		data_out <= r_27_25;
		if (write_en==1'b1)
			r_27_25 <= data_in;
	if (addr_selector[27]&addr_selector[26])
		data_out <= r_27_26;
		if (write_en==1'b1)
			r_27_26 <= data_in;
	if (addr_selector[27]&addr_selector[27])
		data_out <= r_27_27;
		if (write_en==1'b1)
			r_27_27 <= data_in;
	if (addr_selector[27]&addr_selector[28])
		data_out <= r_27_28;
		if (write_en==1'b1)
			r_27_28 <= data_in;
	if (addr_selector[27]&addr_selector[29])
		data_out <= r_27_29;
		if (write_en==1'b1)
			r_27_29 <= data_in;
	if (addr_selector[27]&addr_selector[30])
		data_out <= r_27_30;
		if (write_en==1'b1)
			r_27_30 <= data_in;
	if (addr_selector[27]&addr_selector[31])
		data_out <= r_27_31;
		if (write_en==1'b1)
			r_27_31 <= data_in;
	if (addr_selector[27]&addr_selector[32])
		data_out <= r_27_32;
		if (write_en==1'b1)
			r_27_32 <= data_in;
	if (addr_selector[27]&addr_selector[33])
		data_out <= r_27_33;
		if (write_en==1'b1)
			r_27_33 <= data_in;
	if (addr_selector[27]&addr_selector[34])
		data_out <= r_27_34;
		if (write_en==1'b1)
			r_27_34 <= data_in;
	if (addr_selector[27]&addr_selector[35])
		data_out <= r_27_35;
		if (write_en==1'b1)
			r_27_35 <= data_in;
	if (addr_selector[27]&addr_selector[36])
		data_out <= r_27_36;
		if (write_en==1'b1)
			r_27_36 <= data_in;
	if (addr_selector[27]&addr_selector[37])
		data_out <= r_27_37;
		if (write_en==1'b1)
			r_27_37 <= data_in;
	if (addr_selector[27]&addr_selector[38])
		data_out <= r_27_38;
		if (write_en==1'b1)
			r_27_38 <= data_in;
	if (addr_selector[27]&addr_selector[39])
		data_out <= r_27_39;
		if (write_en==1'b1)
			r_27_39 <= data_in;
	if (addr_selector[27]&addr_selector[40])
		data_out <= r_27_40;
		if (write_en==1'b1)
			r_27_40 <= data_in;
	if (addr_selector[27]&addr_selector[41])
		data_out <= r_27_41;
		if (write_en==1'b1)
			r_27_41 <= data_in;
	if (addr_selector[27]&addr_selector[42])
		data_out <= r_27_42;
		if (write_en==1'b1)
			r_27_42 <= data_in;
	if (addr_selector[27]&addr_selector[43])
		data_out <= r_27_43;
		if (write_en==1'b1)
			r_27_43 <= data_in;
	if (addr_selector[27]&addr_selector[44])
		data_out <= r_27_44;
		if (write_en==1'b1)
			r_27_44 <= data_in;
	if (addr_selector[27]&addr_selector[45])
		data_out <= r_27_45;
		if (write_en==1'b1)
			r_27_45 <= data_in;
	if (addr_selector[27]&addr_selector[46])
		data_out <= r_27_46;
		if (write_en==1'b1)
			r_27_46 <= data_in;
	if (addr_selector[27]&addr_selector[47])
		data_out <= r_27_47;
		if (write_en==1'b1)
			r_27_47 <= data_in;
	if (addr_selector[27]&addr_selector[48])
		data_out <= r_27_48;
		if (write_en==1'b1)
			r_27_48 <= data_in;
	if (addr_selector[27]&addr_selector[49])
		data_out <= r_27_49;
		if (write_en==1'b1)
			r_27_49 <= data_in;
	if (addr_selector[27]&addr_selector[50])
		data_out <= r_27_50;
		if (write_en==1'b1)
			r_27_50 <= data_in;
	if (addr_selector[27]&addr_selector[51])
		data_out <= r_27_51;
		if (write_en==1'b1)
			r_27_51 <= data_in;
	if (addr_selector[27]&addr_selector[52])
		data_out <= r_27_52;
		if (write_en==1'b1)
			r_27_52 <= data_in;
	if (addr_selector[27]&addr_selector[53])
		data_out <= r_27_53;
		if (write_en==1'b1)
			r_27_53 <= data_in;
	if (addr_selector[27]&addr_selector[54])
		data_out <= r_27_54;
		if (write_en==1'b1)
			r_27_54 <= data_in;
	if (addr_selector[27]&addr_selector[55])
		data_out <= r_27_55;
		if (write_en==1'b1)
			r_27_55 <= data_in;
	if (addr_selector[27]&addr_selector[56])
		data_out <= r_27_56;
		if (write_en==1'b1)
			r_27_56 <= data_in;
	if (addr_selector[27]&addr_selector[57])
		data_out <= r_27_57;
		if (write_en==1'b1)
			r_27_57 <= data_in;
	if (addr_selector[27]&addr_selector[58])
		data_out <= r_27_58;
		if (write_en==1'b1)
			r_27_58 <= data_in;
	if (addr_selector[27]&addr_selector[59])
		data_out <= r_27_59;
		if (write_en==1'b1)
			r_27_59 <= data_in;
	if (addr_selector[27]&addr_selector[60])
		data_out <= r_27_60;
		if (write_en==1'b1)
			r_27_60 <= data_in;
	if (addr_selector[27]&addr_selector[61])
		data_out <= r_27_61;
		if (write_en==1'b1)
			r_27_61 <= data_in;
	if (addr_selector[27]&addr_selector[62])
		data_out <= r_27_62;
		if (write_en==1'b1)
			r_27_62 <= data_in;
	if (addr_selector[27]&addr_selector[63])
		data_out <= r_27_63;
		if (write_en==1'b1)
			r_27_63 <= data_in;
	if (addr_selector[28]&addr_selector[0])
		data_out <= r_28_0;
		if (write_en==1'b1)
			r_28_0 <= data_in;
	if (addr_selector[28]&addr_selector[1])
		data_out <= r_28_1;
		if (write_en==1'b1)
			r_28_1 <= data_in;
	if (addr_selector[28]&addr_selector[2])
		data_out <= r_28_2;
		if (write_en==1'b1)
			r_28_2 <= data_in;
	if (addr_selector[28]&addr_selector[3])
		data_out <= r_28_3;
		if (write_en==1'b1)
			r_28_3 <= data_in;
	if (addr_selector[28]&addr_selector[4])
		data_out <= r_28_4;
		if (write_en==1'b1)
			r_28_4 <= data_in;
	if (addr_selector[28]&addr_selector[5])
		data_out <= r_28_5;
		if (write_en==1'b1)
			r_28_5 <= data_in;
	if (addr_selector[28]&addr_selector[6])
		data_out <= r_28_6;
		if (write_en==1'b1)
			r_28_6 <= data_in;
	if (addr_selector[28]&addr_selector[7])
		data_out <= r_28_7;
		if (write_en==1'b1)
			r_28_7 <= data_in;
	if (addr_selector[28]&addr_selector[8])
		data_out <= r_28_8;
		if (write_en==1'b1)
			r_28_8 <= data_in;
	if (addr_selector[28]&addr_selector[9])
		data_out <= r_28_9;
		if (write_en==1'b1)
			r_28_9 <= data_in;
	if (addr_selector[28]&addr_selector[10])
		data_out <= r_28_10;
		if (write_en==1'b1)
			r_28_10 <= data_in;
	if (addr_selector[28]&addr_selector[11])
		data_out <= r_28_11;
		if (write_en==1'b1)
			r_28_11 <= data_in;
	if (addr_selector[28]&addr_selector[12])
		data_out <= r_28_12;
		if (write_en==1'b1)
			r_28_12 <= data_in;
	if (addr_selector[28]&addr_selector[13])
		data_out <= r_28_13;
		if (write_en==1'b1)
			r_28_13 <= data_in;
	if (addr_selector[28]&addr_selector[14])
		data_out <= r_28_14;
		if (write_en==1'b1)
			r_28_14 <= data_in;
	if (addr_selector[28]&addr_selector[15])
		data_out <= r_28_15;
		if (write_en==1'b1)
			r_28_15 <= data_in;
	if (addr_selector[28]&addr_selector[16])
		data_out <= r_28_16;
		if (write_en==1'b1)
			r_28_16 <= data_in;
	if (addr_selector[28]&addr_selector[17])
		data_out <= r_28_17;
		if (write_en==1'b1)
			r_28_17 <= data_in;
	if (addr_selector[28]&addr_selector[18])
		data_out <= r_28_18;
		if (write_en==1'b1)
			r_28_18 <= data_in;
	if (addr_selector[28]&addr_selector[19])
		data_out <= r_28_19;
		if (write_en==1'b1)
			r_28_19 <= data_in;
	if (addr_selector[28]&addr_selector[20])
		data_out <= r_28_20;
		if (write_en==1'b1)
			r_28_20 <= data_in;
	if (addr_selector[28]&addr_selector[21])
		data_out <= r_28_21;
		if (write_en==1'b1)
			r_28_21 <= data_in;
	if (addr_selector[28]&addr_selector[22])
		data_out <= r_28_22;
		if (write_en==1'b1)
			r_28_22 <= data_in;
	if (addr_selector[28]&addr_selector[23])
		data_out <= r_28_23;
		if (write_en==1'b1)
			r_28_23 <= data_in;
	if (addr_selector[28]&addr_selector[24])
		data_out <= r_28_24;
		if (write_en==1'b1)
			r_28_24 <= data_in;
	if (addr_selector[28]&addr_selector[25])
		data_out <= r_28_25;
		if (write_en==1'b1)
			r_28_25 <= data_in;
	if (addr_selector[28]&addr_selector[26])
		data_out <= r_28_26;
		if (write_en==1'b1)
			r_28_26 <= data_in;
	if (addr_selector[28]&addr_selector[27])
		data_out <= r_28_27;
		if (write_en==1'b1)
			r_28_27 <= data_in;
	if (addr_selector[28]&addr_selector[28])
		data_out <= r_28_28;
		if (write_en==1'b1)
			r_28_28 <= data_in;
	if (addr_selector[28]&addr_selector[29])
		data_out <= r_28_29;
		if (write_en==1'b1)
			r_28_29 <= data_in;
	if (addr_selector[28]&addr_selector[30])
		data_out <= r_28_30;
		if (write_en==1'b1)
			r_28_30 <= data_in;
	if (addr_selector[28]&addr_selector[31])
		data_out <= r_28_31;
		if (write_en==1'b1)
			r_28_31 <= data_in;
	if (addr_selector[28]&addr_selector[32])
		data_out <= r_28_32;
		if (write_en==1'b1)
			r_28_32 <= data_in;
	if (addr_selector[28]&addr_selector[33])
		data_out <= r_28_33;
		if (write_en==1'b1)
			r_28_33 <= data_in;
	if (addr_selector[28]&addr_selector[34])
		data_out <= r_28_34;
		if (write_en==1'b1)
			r_28_34 <= data_in;
	if (addr_selector[28]&addr_selector[35])
		data_out <= r_28_35;
		if (write_en==1'b1)
			r_28_35 <= data_in;
	if (addr_selector[28]&addr_selector[36])
		data_out <= r_28_36;
		if (write_en==1'b1)
			r_28_36 <= data_in;
	if (addr_selector[28]&addr_selector[37])
		data_out <= r_28_37;
		if (write_en==1'b1)
			r_28_37 <= data_in;
	if (addr_selector[28]&addr_selector[38])
		data_out <= r_28_38;
		if (write_en==1'b1)
			r_28_38 <= data_in;
	if (addr_selector[28]&addr_selector[39])
		data_out <= r_28_39;
		if (write_en==1'b1)
			r_28_39 <= data_in;
	if (addr_selector[28]&addr_selector[40])
		data_out <= r_28_40;
		if (write_en==1'b1)
			r_28_40 <= data_in;
	if (addr_selector[28]&addr_selector[41])
		data_out <= r_28_41;
		if (write_en==1'b1)
			r_28_41 <= data_in;
	if (addr_selector[28]&addr_selector[42])
		data_out <= r_28_42;
		if (write_en==1'b1)
			r_28_42 <= data_in;
	if (addr_selector[28]&addr_selector[43])
		data_out <= r_28_43;
		if (write_en==1'b1)
			r_28_43 <= data_in;
	if (addr_selector[28]&addr_selector[44])
		data_out <= r_28_44;
		if (write_en==1'b1)
			r_28_44 <= data_in;
	if (addr_selector[28]&addr_selector[45])
		data_out <= r_28_45;
		if (write_en==1'b1)
			r_28_45 <= data_in;
	if (addr_selector[28]&addr_selector[46])
		data_out <= r_28_46;
		if (write_en==1'b1)
			r_28_46 <= data_in;
	if (addr_selector[28]&addr_selector[47])
		data_out <= r_28_47;
		if (write_en==1'b1)
			r_28_47 <= data_in;
	if (addr_selector[28]&addr_selector[48])
		data_out <= r_28_48;
		if (write_en==1'b1)
			r_28_48 <= data_in;
	if (addr_selector[28]&addr_selector[49])
		data_out <= r_28_49;
		if (write_en==1'b1)
			r_28_49 <= data_in;
	if (addr_selector[28]&addr_selector[50])
		data_out <= r_28_50;
		if (write_en==1'b1)
			r_28_50 <= data_in;
	if (addr_selector[28]&addr_selector[51])
		data_out <= r_28_51;
		if (write_en==1'b1)
			r_28_51 <= data_in;
	if (addr_selector[28]&addr_selector[52])
		data_out <= r_28_52;
		if (write_en==1'b1)
			r_28_52 <= data_in;
	if (addr_selector[28]&addr_selector[53])
		data_out <= r_28_53;
		if (write_en==1'b1)
			r_28_53 <= data_in;
	if (addr_selector[28]&addr_selector[54])
		data_out <= r_28_54;
		if (write_en==1'b1)
			r_28_54 <= data_in;
	if (addr_selector[28]&addr_selector[55])
		data_out <= r_28_55;
		if (write_en==1'b1)
			r_28_55 <= data_in;
	if (addr_selector[28]&addr_selector[56])
		data_out <= r_28_56;
		if (write_en==1'b1)
			r_28_56 <= data_in;
	if (addr_selector[28]&addr_selector[57])
		data_out <= r_28_57;
		if (write_en==1'b1)
			r_28_57 <= data_in;
	if (addr_selector[28]&addr_selector[58])
		data_out <= r_28_58;
		if (write_en==1'b1)
			r_28_58 <= data_in;
	if (addr_selector[28]&addr_selector[59])
		data_out <= r_28_59;
		if (write_en==1'b1)
			r_28_59 <= data_in;
	if (addr_selector[28]&addr_selector[60])
		data_out <= r_28_60;
		if (write_en==1'b1)
			r_28_60 <= data_in;
	if (addr_selector[28]&addr_selector[61])
		data_out <= r_28_61;
		if (write_en==1'b1)
			r_28_61 <= data_in;
	if (addr_selector[28]&addr_selector[62])
		data_out <= r_28_62;
		if (write_en==1'b1)
			r_28_62 <= data_in;
	if (addr_selector[28]&addr_selector[63])
		data_out <= r_28_63;
		if (write_en==1'b1)
			r_28_63 <= data_in;
	if (addr_selector[29]&addr_selector[0])
		data_out <= r_29_0;
		if (write_en==1'b1)
			r_29_0 <= data_in;
	if (addr_selector[29]&addr_selector[1])
		data_out <= r_29_1;
		if (write_en==1'b1)
			r_29_1 <= data_in;
	if (addr_selector[29]&addr_selector[2])
		data_out <= r_29_2;
		if (write_en==1'b1)
			r_29_2 <= data_in;
	if (addr_selector[29]&addr_selector[3])
		data_out <= r_29_3;
		if (write_en==1'b1)
			r_29_3 <= data_in;
	if (addr_selector[29]&addr_selector[4])
		data_out <= r_29_4;
		if (write_en==1'b1)
			r_29_4 <= data_in;
	if (addr_selector[29]&addr_selector[5])
		data_out <= r_29_5;
		if (write_en==1'b1)
			r_29_5 <= data_in;
	if (addr_selector[29]&addr_selector[6])
		data_out <= r_29_6;
		if (write_en==1'b1)
			r_29_6 <= data_in;
	if (addr_selector[29]&addr_selector[7])
		data_out <= r_29_7;
		if (write_en==1'b1)
			r_29_7 <= data_in;
	if (addr_selector[29]&addr_selector[8])
		data_out <= r_29_8;
		if (write_en==1'b1)
			r_29_8 <= data_in;
	if (addr_selector[29]&addr_selector[9])
		data_out <= r_29_9;
		if (write_en==1'b1)
			r_29_9 <= data_in;
	if (addr_selector[29]&addr_selector[10])
		data_out <= r_29_10;
		if (write_en==1'b1)
			r_29_10 <= data_in;
	if (addr_selector[29]&addr_selector[11])
		data_out <= r_29_11;
		if (write_en==1'b1)
			r_29_11 <= data_in;
	if (addr_selector[29]&addr_selector[12])
		data_out <= r_29_12;
		if (write_en==1'b1)
			r_29_12 <= data_in;
	if (addr_selector[29]&addr_selector[13])
		data_out <= r_29_13;
		if (write_en==1'b1)
			r_29_13 <= data_in;
	if (addr_selector[29]&addr_selector[14])
		data_out <= r_29_14;
		if (write_en==1'b1)
			r_29_14 <= data_in;
	if (addr_selector[29]&addr_selector[15])
		data_out <= r_29_15;
		if (write_en==1'b1)
			r_29_15 <= data_in;
	if (addr_selector[29]&addr_selector[16])
		data_out <= r_29_16;
		if (write_en==1'b1)
			r_29_16 <= data_in;
	if (addr_selector[29]&addr_selector[17])
		data_out <= r_29_17;
		if (write_en==1'b1)
			r_29_17 <= data_in;
	if (addr_selector[29]&addr_selector[18])
		data_out <= r_29_18;
		if (write_en==1'b1)
			r_29_18 <= data_in;
	if (addr_selector[29]&addr_selector[19])
		data_out <= r_29_19;
		if (write_en==1'b1)
			r_29_19 <= data_in;
	if (addr_selector[29]&addr_selector[20])
		data_out <= r_29_20;
		if (write_en==1'b1)
			r_29_20 <= data_in;
	if (addr_selector[29]&addr_selector[21])
		data_out <= r_29_21;
		if (write_en==1'b1)
			r_29_21 <= data_in;
	if (addr_selector[29]&addr_selector[22])
		data_out <= r_29_22;
		if (write_en==1'b1)
			r_29_22 <= data_in;
	if (addr_selector[29]&addr_selector[23])
		data_out <= r_29_23;
		if (write_en==1'b1)
			r_29_23 <= data_in;
	if (addr_selector[29]&addr_selector[24])
		data_out <= r_29_24;
		if (write_en==1'b1)
			r_29_24 <= data_in;
	if (addr_selector[29]&addr_selector[25])
		data_out <= r_29_25;
		if (write_en==1'b1)
			r_29_25 <= data_in;
	if (addr_selector[29]&addr_selector[26])
		data_out <= r_29_26;
		if (write_en==1'b1)
			r_29_26 <= data_in;
	if (addr_selector[29]&addr_selector[27])
		data_out <= r_29_27;
		if (write_en==1'b1)
			r_29_27 <= data_in;
	if (addr_selector[29]&addr_selector[28])
		data_out <= r_29_28;
		if (write_en==1'b1)
			r_29_28 <= data_in;
	if (addr_selector[29]&addr_selector[29])
		data_out <= r_29_29;
		if (write_en==1'b1)
			r_29_29 <= data_in;
	if (addr_selector[29]&addr_selector[30])
		data_out <= r_29_30;
		if (write_en==1'b1)
			r_29_30 <= data_in;
	if (addr_selector[29]&addr_selector[31])
		data_out <= r_29_31;
		if (write_en==1'b1)
			r_29_31 <= data_in;
	if (addr_selector[29]&addr_selector[32])
		data_out <= r_29_32;
		if (write_en==1'b1)
			r_29_32 <= data_in;
	if (addr_selector[29]&addr_selector[33])
		data_out <= r_29_33;
		if (write_en==1'b1)
			r_29_33 <= data_in;
	if (addr_selector[29]&addr_selector[34])
		data_out <= r_29_34;
		if (write_en==1'b1)
			r_29_34 <= data_in;
	if (addr_selector[29]&addr_selector[35])
		data_out <= r_29_35;
		if (write_en==1'b1)
			r_29_35 <= data_in;
	if (addr_selector[29]&addr_selector[36])
		data_out <= r_29_36;
		if (write_en==1'b1)
			r_29_36 <= data_in;
	if (addr_selector[29]&addr_selector[37])
		data_out <= r_29_37;
		if (write_en==1'b1)
			r_29_37 <= data_in;
	if (addr_selector[29]&addr_selector[38])
		data_out <= r_29_38;
		if (write_en==1'b1)
			r_29_38 <= data_in;
	if (addr_selector[29]&addr_selector[39])
		data_out <= r_29_39;
		if (write_en==1'b1)
			r_29_39 <= data_in;
	if (addr_selector[29]&addr_selector[40])
		data_out <= r_29_40;
		if (write_en==1'b1)
			r_29_40 <= data_in;
	if (addr_selector[29]&addr_selector[41])
		data_out <= r_29_41;
		if (write_en==1'b1)
			r_29_41 <= data_in;
	if (addr_selector[29]&addr_selector[42])
		data_out <= r_29_42;
		if (write_en==1'b1)
			r_29_42 <= data_in;
	if (addr_selector[29]&addr_selector[43])
		data_out <= r_29_43;
		if (write_en==1'b1)
			r_29_43 <= data_in;
	if (addr_selector[29]&addr_selector[44])
		data_out <= r_29_44;
		if (write_en==1'b1)
			r_29_44 <= data_in;
	if (addr_selector[29]&addr_selector[45])
		data_out <= r_29_45;
		if (write_en==1'b1)
			r_29_45 <= data_in;
	if (addr_selector[29]&addr_selector[46])
		data_out <= r_29_46;
		if (write_en==1'b1)
			r_29_46 <= data_in;
	if (addr_selector[29]&addr_selector[47])
		data_out <= r_29_47;
		if (write_en==1'b1)
			r_29_47 <= data_in;
	if (addr_selector[29]&addr_selector[48])
		data_out <= r_29_48;
		if (write_en==1'b1)
			r_29_48 <= data_in;
	if (addr_selector[29]&addr_selector[49])
		data_out <= r_29_49;
		if (write_en==1'b1)
			r_29_49 <= data_in;
	if (addr_selector[29]&addr_selector[50])
		data_out <= r_29_50;
		if (write_en==1'b1)
			r_29_50 <= data_in;
	if (addr_selector[29]&addr_selector[51])
		data_out <= r_29_51;
		if (write_en==1'b1)
			r_29_51 <= data_in;
	if (addr_selector[29]&addr_selector[52])
		data_out <= r_29_52;
		if (write_en==1'b1)
			r_29_52 <= data_in;
	if (addr_selector[29]&addr_selector[53])
		data_out <= r_29_53;
		if (write_en==1'b1)
			r_29_53 <= data_in;
	if (addr_selector[29]&addr_selector[54])
		data_out <= r_29_54;
		if (write_en==1'b1)
			r_29_54 <= data_in;
	if (addr_selector[29]&addr_selector[55])
		data_out <= r_29_55;
		if (write_en==1'b1)
			r_29_55 <= data_in;
	if (addr_selector[29]&addr_selector[56])
		data_out <= r_29_56;
		if (write_en==1'b1)
			r_29_56 <= data_in;
	if (addr_selector[29]&addr_selector[57])
		data_out <= r_29_57;
		if (write_en==1'b1)
			r_29_57 <= data_in;
	if (addr_selector[29]&addr_selector[58])
		data_out <= r_29_58;
		if (write_en==1'b1)
			r_29_58 <= data_in;
	if (addr_selector[29]&addr_selector[59])
		data_out <= r_29_59;
		if (write_en==1'b1)
			r_29_59 <= data_in;
	if (addr_selector[29]&addr_selector[60])
		data_out <= r_29_60;
		if (write_en==1'b1)
			r_29_60 <= data_in;
	if (addr_selector[29]&addr_selector[61])
		data_out <= r_29_61;
		if (write_en==1'b1)
			r_29_61 <= data_in;
	if (addr_selector[29]&addr_selector[62])
		data_out <= r_29_62;
		if (write_en==1'b1)
			r_29_62 <= data_in;
	if (addr_selector[29]&addr_selector[63])
		data_out <= r_29_63;
		if (write_en==1'b1)
			r_29_63 <= data_in;
	if (addr_selector[30]&addr_selector[0])
		data_out <= r_30_0;
		if (write_en==1'b1)
			r_30_0 <= data_in;
	if (addr_selector[30]&addr_selector[1])
		data_out <= r_30_1;
		if (write_en==1'b1)
			r_30_1 <= data_in;
	if (addr_selector[30]&addr_selector[2])
		data_out <= r_30_2;
		if (write_en==1'b1)
			r_30_2 <= data_in;
	if (addr_selector[30]&addr_selector[3])
		data_out <= r_30_3;
		if (write_en==1'b1)
			r_30_3 <= data_in;
	if (addr_selector[30]&addr_selector[4])
		data_out <= r_30_4;
		if (write_en==1'b1)
			r_30_4 <= data_in;
	if (addr_selector[30]&addr_selector[5])
		data_out <= r_30_5;
		if (write_en==1'b1)
			r_30_5 <= data_in;
	if (addr_selector[30]&addr_selector[6])
		data_out <= r_30_6;
		if (write_en==1'b1)
			r_30_6 <= data_in;
	if (addr_selector[30]&addr_selector[7])
		data_out <= r_30_7;
		if (write_en==1'b1)
			r_30_7 <= data_in;
	if (addr_selector[30]&addr_selector[8])
		data_out <= r_30_8;
		if (write_en==1'b1)
			r_30_8 <= data_in;
	if (addr_selector[30]&addr_selector[9])
		data_out <= r_30_9;
		if (write_en==1'b1)
			r_30_9 <= data_in;
	if (addr_selector[30]&addr_selector[10])
		data_out <= r_30_10;
		if (write_en==1'b1)
			r_30_10 <= data_in;
	if (addr_selector[30]&addr_selector[11])
		data_out <= r_30_11;
		if (write_en==1'b1)
			r_30_11 <= data_in;
	if (addr_selector[30]&addr_selector[12])
		data_out <= r_30_12;
		if (write_en==1'b1)
			r_30_12 <= data_in;
	if (addr_selector[30]&addr_selector[13])
		data_out <= r_30_13;
		if (write_en==1'b1)
			r_30_13 <= data_in;
	if (addr_selector[30]&addr_selector[14])
		data_out <= r_30_14;
		if (write_en==1'b1)
			r_30_14 <= data_in;
	if (addr_selector[30]&addr_selector[15])
		data_out <= r_30_15;
		if (write_en==1'b1)
			r_30_15 <= data_in;
	if (addr_selector[30]&addr_selector[16])
		data_out <= r_30_16;
		if (write_en==1'b1)
			r_30_16 <= data_in;
	if (addr_selector[30]&addr_selector[17])
		data_out <= r_30_17;
		if (write_en==1'b1)
			r_30_17 <= data_in;
	if (addr_selector[30]&addr_selector[18])
		data_out <= r_30_18;
		if (write_en==1'b1)
			r_30_18 <= data_in;
	if (addr_selector[30]&addr_selector[19])
		data_out <= r_30_19;
		if (write_en==1'b1)
			r_30_19 <= data_in;
	if (addr_selector[30]&addr_selector[20])
		data_out <= r_30_20;
		if (write_en==1'b1)
			r_30_20 <= data_in;
	if (addr_selector[30]&addr_selector[21])
		data_out <= r_30_21;
		if (write_en==1'b1)
			r_30_21 <= data_in;
	if (addr_selector[30]&addr_selector[22])
		data_out <= r_30_22;
		if (write_en==1'b1)
			r_30_22 <= data_in;
	if (addr_selector[30]&addr_selector[23])
		data_out <= r_30_23;
		if (write_en==1'b1)
			r_30_23 <= data_in;
	if (addr_selector[30]&addr_selector[24])
		data_out <= r_30_24;
		if (write_en==1'b1)
			r_30_24 <= data_in;
	if (addr_selector[30]&addr_selector[25])
		data_out <= r_30_25;
		if (write_en==1'b1)
			r_30_25 <= data_in;
	if (addr_selector[30]&addr_selector[26])
		data_out <= r_30_26;
		if (write_en==1'b1)
			r_30_26 <= data_in;
	if (addr_selector[30]&addr_selector[27])
		data_out <= r_30_27;
		if (write_en==1'b1)
			r_30_27 <= data_in;
	if (addr_selector[30]&addr_selector[28])
		data_out <= r_30_28;
		if (write_en==1'b1)
			r_30_28 <= data_in;
	if (addr_selector[30]&addr_selector[29])
		data_out <= r_30_29;
		if (write_en==1'b1)
			r_30_29 <= data_in;
	if (addr_selector[30]&addr_selector[30])
		data_out <= r_30_30;
		if (write_en==1'b1)
			r_30_30 <= data_in;
	if (addr_selector[30]&addr_selector[31])
		data_out <= r_30_31;
		if (write_en==1'b1)
			r_30_31 <= data_in;
	if (addr_selector[30]&addr_selector[32])
		data_out <= r_30_32;
		if (write_en==1'b1)
			r_30_32 <= data_in;
	if (addr_selector[30]&addr_selector[33])
		data_out <= r_30_33;
		if (write_en==1'b1)
			r_30_33 <= data_in;
	if (addr_selector[30]&addr_selector[34])
		data_out <= r_30_34;
		if (write_en==1'b1)
			r_30_34 <= data_in;
	if (addr_selector[30]&addr_selector[35])
		data_out <= r_30_35;
		if (write_en==1'b1)
			r_30_35 <= data_in;
	if (addr_selector[30]&addr_selector[36])
		data_out <= r_30_36;
		if (write_en==1'b1)
			r_30_36 <= data_in;
	if (addr_selector[30]&addr_selector[37])
		data_out <= r_30_37;
		if (write_en==1'b1)
			r_30_37 <= data_in;
	if (addr_selector[30]&addr_selector[38])
		data_out <= r_30_38;
		if (write_en==1'b1)
			r_30_38 <= data_in;
	if (addr_selector[30]&addr_selector[39])
		data_out <= r_30_39;
		if (write_en==1'b1)
			r_30_39 <= data_in;
	if (addr_selector[30]&addr_selector[40])
		data_out <= r_30_40;
		if (write_en==1'b1)
			r_30_40 <= data_in;
	if (addr_selector[30]&addr_selector[41])
		data_out <= r_30_41;
		if (write_en==1'b1)
			r_30_41 <= data_in;
	if (addr_selector[30]&addr_selector[42])
		data_out <= r_30_42;
		if (write_en==1'b1)
			r_30_42 <= data_in;
	if (addr_selector[30]&addr_selector[43])
		data_out <= r_30_43;
		if (write_en==1'b1)
			r_30_43 <= data_in;
	if (addr_selector[30]&addr_selector[44])
		data_out <= r_30_44;
		if (write_en==1'b1)
			r_30_44 <= data_in;
	if (addr_selector[30]&addr_selector[45])
		data_out <= r_30_45;
		if (write_en==1'b1)
			r_30_45 <= data_in;
	if (addr_selector[30]&addr_selector[46])
		data_out <= r_30_46;
		if (write_en==1'b1)
			r_30_46 <= data_in;
	if (addr_selector[30]&addr_selector[47])
		data_out <= r_30_47;
		if (write_en==1'b1)
			r_30_47 <= data_in;
	if (addr_selector[30]&addr_selector[48])
		data_out <= r_30_48;
		if (write_en==1'b1)
			r_30_48 <= data_in;
	if (addr_selector[30]&addr_selector[49])
		data_out <= r_30_49;
		if (write_en==1'b1)
			r_30_49 <= data_in;
	if (addr_selector[30]&addr_selector[50])
		data_out <= r_30_50;
		if (write_en==1'b1)
			r_30_50 <= data_in;
	if (addr_selector[30]&addr_selector[51])
		data_out <= r_30_51;
		if (write_en==1'b1)
			r_30_51 <= data_in;
	if (addr_selector[30]&addr_selector[52])
		data_out <= r_30_52;
		if (write_en==1'b1)
			r_30_52 <= data_in;
	if (addr_selector[30]&addr_selector[53])
		data_out <= r_30_53;
		if (write_en==1'b1)
			r_30_53 <= data_in;
	if (addr_selector[30]&addr_selector[54])
		data_out <= r_30_54;
		if (write_en==1'b1)
			r_30_54 <= data_in;
	if (addr_selector[30]&addr_selector[55])
		data_out <= r_30_55;
		if (write_en==1'b1)
			r_30_55 <= data_in;
	if (addr_selector[30]&addr_selector[56])
		data_out <= r_30_56;
		if (write_en==1'b1)
			r_30_56 <= data_in;
	if (addr_selector[30]&addr_selector[57])
		data_out <= r_30_57;
		if (write_en==1'b1)
			r_30_57 <= data_in;
	if (addr_selector[30]&addr_selector[58])
		data_out <= r_30_58;
		if (write_en==1'b1)
			r_30_58 <= data_in;
	if (addr_selector[30]&addr_selector[59])
		data_out <= r_30_59;
		if (write_en==1'b1)
			r_30_59 <= data_in;
	if (addr_selector[30]&addr_selector[60])
		data_out <= r_30_60;
		if (write_en==1'b1)
			r_30_60 <= data_in;
	if (addr_selector[30]&addr_selector[61])
		data_out <= r_30_61;
		if (write_en==1'b1)
			r_30_61 <= data_in;
	if (addr_selector[30]&addr_selector[62])
		data_out <= r_30_62;
		if (write_en==1'b1)
			r_30_62 <= data_in;
	if (addr_selector[30]&addr_selector[63])
		data_out <= r_30_63;
		if (write_en==1'b1)
			r_30_63 <= data_in;
	if (addr_selector[31]&addr_selector[0])
		data_out <= r_31_0;
		if (write_en==1'b1)
			r_31_0 <= data_in;
	if (addr_selector[31]&addr_selector[1])
		data_out <= r_31_1;
		if (write_en==1'b1)
			r_31_1 <= data_in;
	if (addr_selector[31]&addr_selector[2])
		data_out <= r_31_2;
		if (write_en==1'b1)
			r_31_2 <= data_in;
	if (addr_selector[31]&addr_selector[3])
		data_out <= r_31_3;
		if (write_en==1'b1)
			r_31_3 <= data_in;
	if (addr_selector[31]&addr_selector[4])
		data_out <= r_31_4;
		if (write_en==1'b1)
			r_31_4 <= data_in;
	if (addr_selector[31]&addr_selector[5])
		data_out <= r_31_5;
		if (write_en==1'b1)
			r_31_5 <= data_in;
	if (addr_selector[31]&addr_selector[6])
		data_out <= r_31_6;
		if (write_en==1'b1)
			r_31_6 <= data_in;
	if (addr_selector[31]&addr_selector[7])
		data_out <= r_31_7;
		if (write_en==1'b1)
			r_31_7 <= data_in;
	if (addr_selector[31]&addr_selector[8])
		data_out <= r_31_8;
		if (write_en==1'b1)
			r_31_8 <= data_in;
	if (addr_selector[31]&addr_selector[9])
		data_out <= r_31_9;
		if (write_en==1'b1)
			r_31_9 <= data_in;
	if (addr_selector[31]&addr_selector[10])
		data_out <= r_31_10;
		if (write_en==1'b1)
			r_31_10 <= data_in;
	if (addr_selector[31]&addr_selector[11])
		data_out <= r_31_11;
		if (write_en==1'b1)
			r_31_11 <= data_in;
	if (addr_selector[31]&addr_selector[12])
		data_out <= r_31_12;
		if (write_en==1'b1)
			r_31_12 <= data_in;
	if (addr_selector[31]&addr_selector[13])
		data_out <= r_31_13;
		if (write_en==1'b1)
			r_31_13 <= data_in;
	if (addr_selector[31]&addr_selector[14])
		data_out <= r_31_14;
		if (write_en==1'b1)
			r_31_14 <= data_in;
	if (addr_selector[31]&addr_selector[15])
		data_out <= r_31_15;
		if (write_en==1'b1)
			r_31_15 <= data_in;
	if (addr_selector[31]&addr_selector[16])
		data_out <= r_31_16;
		if (write_en==1'b1)
			r_31_16 <= data_in;
	if (addr_selector[31]&addr_selector[17])
		data_out <= r_31_17;
		if (write_en==1'b1)
			r_31_17 <= data_in;
	if (addr_selector[31]&addr_selector[18])
		data_out <= r_31_18;
		if (write_en==1'b1)
			r_31_18 <= data_in;
	if (addr_selector[31]&addr_selector[19])
		data_out <= r_31_19;
		if (write_en==1'b1)
			r_31_19 <= data_in;
	if (addr_selector[31]&addr_selector[20])
		data_out <= r_31_20;
		if (write_en==1'b1)
			r_31_20 <= data_in;
	if (addr_selector[31]&addr_selector[21])
		data_out <= r_31_21;
		if (write_en==1'b1)
			r_31_21 <= data_in;
	if (addr_selector[31]&addr_selector[22])
		data_out <= r_31_22;
		if (write_en==1'b1)
			r_31_22 <= data_in;
	if (addr_selector[31]&addr_selector[23])
		data_out <= r_31_23;
		if (write_en==1'b1)
			r_31_23 <= data_in;
	if (addr_selector[31]&addr_selector[24])
		data_out <= r_31_24;
		if (write_en==1'b1)
			r_31_24 <= data_in;
	if (addr_selector[31]&addr_selector[25])
		data_out <= r_31_25;
		if (write_en==1'b1)
			r_31_25 <= data_in;
	if (addr_selector[31]&addr_selector[26])
		data_out <= r_31_26;
		if (write_en==1'b1)
			r_31_26 <= data_in;
	if (addr_selector[31]&addr_selector[27])
		data_out <= r_31_27;
		if (write_en==1'b1)
			r_31_27 <= data_in;
	if (addr_selector[31]&addr_selector[28])
		data_out <= r_31_28;
		if (write_en==1'b1)
			r_31_28 <= data_in;
	if (addr_selector[31]&addr_selector[29])
		data_out <= r_31_29;
		if (write_en==1'b1)
			r_31_29 <= data_in;
	if (addr_selector[31]&addr_selector[30])
		data_out <= r_31_30;
		if (write_en==1'b1)
			r_31_30 <= data_in;
	if (addr_selector[31]&addr_selector[31])
		data_out <= r_31_31;
		if (write_en==1'b1)
			r_31_31 <= data_in;
	if (addr_selector[31]&addr_selector[32])
		data_out <= r_31_32;
		if (write_en==1'b1)
			r_31_32 <= data_in;
	if (addr_selector[31]&addr_selector[33])
		data_out <= r_31_33;
		if (write_en==1'b1)
			r_31_33 <= data_in;
	if (addr_selector[31]&addr_selector[34])
		data_out <= r_31_34;
		if (write_en==1'b1)
			r_31_34 <= data_in;
	if (addr_selector[31]&addr_selector[35])
		data_out <= r_31_35;
		if (write_en==1'b1)
			r_31_35 <= data_in;
	if (addr_selector[31]&addr_selector[36])
		data_out <= r_31_36;
		if (write_en==1'b1)
			r_31_36 <= data_in;
	if (addr_selector[31]&addr_selector[37])
		data_out <= r_31_37;
		if (write_en==1'b1)
			r_31_37 <= data_in;
	if (addr_selector[31]&addr_selector[38])
		data_out <= r_31_38;
		if (write_en==1'b1)
			r_31_38 <= data_in;
	if (addr_selector[31]&addr_selector[39])
		data_out <= r_31_39;
		if (write_en==1'b1)
			r_31_39 <= data_in;
	if (addr_selector[31]&addr_selector[40])
		data_out <= r_31_40;
		if (write_en==1'b1)
			r_31_40 <= data_in;
	if (addr_selector[31]&addr_selector[41])
		data_out <= r_31_41;
		if (write_en==1'b1)
			r_31_41 <= data_in;
	if (addr_selector[31]&addr_selector[42])
		data_out <= r_31_42;
		if (write_en==1'b1)
			r_31_42 <= data_in;
	if (addr_selector[31]&addr_selector[43])
		data_out <= r_31_43;
		if (write_en==1'b1)
			r_31_43 <= data_in;
	if (addr_selector[31]&addr_selector[44])
		data_out <= r_31_44;
		if (write_en==1'b1)
			r_31_44 <= data_in;
	if (addr_selector[31]&addr_selector[45])
		data_out <= r_31_45;
		if (write_en==1'b1)
			r_31_45 <= data_in;
	if (addr_selector[31]&addr_selector[46])
		data_out <= r_31_46;
		if (write_en==1'b1)
			r_31_46 <= data_in;
	if (addr_selector[31]&addr_selector[47])
		data_out <= r_31_47;
		if (write_en==1'b1)
			r_31_47 <= data_in;
	if (addr_selector[31]&addr_selector[48])
		data_out <= r_31_48;
		if (write_en==1'b1)
			r_31_48 <= data_in;
	if (addr_selector[31]&addr_selector[49])
		data_out <= r_31_49;
		if (write_en==1'b1)
			r_31_49 <= data_in;
	if (addr_selector[31]&addr_selector[50])
		data_out <= r_31_50;
		if (write_en==1'b1)
			r_31_50 <= data_in;
	if (addr_selector[31]&addr_selector[51])
		data_out <= r_31_51;
		if (write_en==1'b1)
			r_31_51 <= data_in;
	if (addr_selector[31]&addr_selector[52])
		data_out <= r_31_52;
		if (write_en==1'b1)
			r_31_52 <= data_in;
	if (addr_selector[31]&addr_selector[53])
		data_out <= r_31_53;
		if (write_en==1'b1)
			r_31_53 <= data_in;
	if (addr_selector[31]&addr_selector[54])
		data_out <= r_31_54;
		if (write_en==1'b1)
			r_31_54 <= data_in;
	if (addr_selector[31]&addr_selector[55])
		data_out <= r_31_55;
		if (write_en==1'b1)
			r_31_55 <= data_in;
	if (addr_selector[31]&addr_selector[56])
		data_out <= r_31_56;
		if (write_en==1'b1)
			r_31_56 <= data_in;
	if (addr_selector[31]&addr_selector[57])
		data_out <= r_31_57;
		if (write_en==1'b1)
			r_31_57 <= data_in;
	if (addr_selector[31]&addr_selector[58])
		data_out <= r_31_58;
		if (write_en==1'b1)
			r_31_58 <= data_in;
	if (addr_selector[31]&addr_selector[59])
		data_out <= r_31_59;
		if (write_en==1'b1)
			r_31_59 <= data_in;
	if (addr_selector[31]&addr_selector[60])
		data_out <= r_31_60;
		if (write_en==1'b1)
			r_31_60 <= data_in;
	if (addr_selector[31]&addr_selector[61])
		data_out <= r_31_61;
		if (write_en==1'b1)
			r_31_61 <= data_in;
	if (addr_selector[31]&addr_selector[62])
		data_out <= r_31_62;
		if (write_en==1'b1)
			r_31_62 <= data_in;
	if (addr_selector[31]&addr_selector[63])
		data_out <= r_31_63;
		if (write_en==1'b1)
			r_31_63 <= data_in;
	if (addr_selector[32]&addr_selector[0])
		data_out <= r_32_0;
		if (write_en==1'b1)
			r_32_0 <= data_in;
	if (addr_selector[32]&addr_selector[1])
		data_out <= r_32_1;
		if (write_en==1'b1)
			r_32_1 <= data_in;
	if (addr_selector[32]&addr_selector[2])
		data_out <= r_32_2;
		if (write_en==1'b1)
			r_32_2 <= data_in;
	if (addr_selector[32]&addr_selector[3])
		data_out <= r_32_3;
		if (write_en==1'b1)
			r_32_3 <= data_in;
	if (addr_selector[32]&addr_selector[4])
		data_out <= r_32_4;
		if (write_en==1'b1)
			r_32_4 <= data_in;
	if (addr_selector[32]&addr_selector[5])
		data_out <= r_32_5;
		if (write_en==1'b1)
			r_32_5 <= data_in;
	if (addr_selector[32]&addr_selector[6])
		data_out <= r_32_6;
		if (write_en==1'b1)
			r_32_6 <= data_in;
	if (addr_selector[32]&addr_selector[7])
		data_out <= r_32_7;
		if (write_en==1'b1)
			r_32_7 <= data_in;
	if (addr_selector[32]&addr_selector[8])
		data_out <= r_32_8;
		if (write_en==1'b1)
			r_32_8 <= data_in;
	if (addr_selector[32]&addr_selector[9])
		data_out <= r_32_9;
		if (write_en==1'b1)
			r_32_9 <= data_in;
	if (addr_selector[32]&addr_selector[10])
		data_out <= r_32_10;
		if (write_en==1'b1)
			r_32_10 <= data_in;
	if (addr_selector[32]&addr_selector[11])
		data_out <= r_32_11;
		if (write_en==1'b1)
			r_32_11 <= data_in;
	if (addr_selector[32]&addr_selector[12])
		data_out <= r_32_12;
		if (write_en==1'b1)
			r_32_12 <= data_in;
	if (addr_selector[32]&addr_selector[13])
		data_out <= r_32_13;
		if (write_en==1'b1)
			r_32_13 <= data_in;
	if (addr_selector[32]&addr_selector[14])
		data_out <= r_32_14;
		if (write_en==1'b1)
			r_32_14 <= data_in;
	if (addr_selector[32]&addr_selector[15])
		data_out <= r_32_15;
		if (write_en==1'b1)
			r_32_15 <= data_in;
	if (addr_selector[32]&addr_selector[16])
		data_out <= r_32_16;
		if (write_en==1'b1)
			r_32_16 <= data_in;
	if (addr_selector[32]&addr_selector[17])
		data_out <= r_32_17;
		if (write_en==1'b1)
			r_32_17 <= data_in;
	if (addr_selector[32]&addr_selector[18])
		data_out <= r_32_18;
		if (write_en==1'b1)
			r_32_18 <= data_in;
	if (addr_selector[32]&addr_selector[19])
		data_out <= r_32_19;
		if (write_en==1'b1)
			r_32_19 <= data_in;
	if (addr_selector[32]&addr_selector[20])
		data_out <= r_32_20;
		if (write_en==1'b1)
			r_32_20 <= data_in;
	if (addr_selector[32]&addr_selector[21])
		data_out <= r_32_21;
		if (write_en==1'b1)
			r_32_21 <= data_in;
	if (addr_selector[32]&addr_selector[22])
		data_out <= r_32_22;
		if (write_en==1'b1)
			r_32_22 <= data_in;
	if (addr_selector[32]&addr_selector[23])
		data_out <= r_32_23;
		if (write_en==1'b1)
			r_32_23 <= data_in;
	if (addr_selector[32]&addr_selector[24])
		data_out <= r_32_24;
		if (write_en==1'b1)
			r_32_24 <= data_in;
	if (addr_selector[32]&addr_selector[25])
		data_out <= r_32_25;
		if (write_en==1'b1)
			r_32_25 <= data_in;
	if (addr_selector[32]&addr_selector[26])
		data_out <= r_32_26;
		if (write_en==1'b1)
			r_32_26 <= data_in;
	if (addr_selector[32]&addr_selector[27])
		data_out <= r_32_27;
		if (write_en==1'b1)
			r_32_27 <= data_in;
	if (addr_selector[32]&addr_selector[28])
		data_out <= r_32_28;
		if (write_en==1'b1)
			r_32_28 <= data_in;
	if (addr_selector[32]&addr_selector[29])
		data_out <= r_32_29;
		if (write_en==1'b1)
			r_32_29 <= data_in;
	if (addr_selector[32]&addr_selector[30])
		data_out <= r_32_30;
		if (write_en==1'b1)
			r_32_30 <= data_in;
	if (addr_selector[32]&addr_selector[31])
		data_out <= r_32_31;
		if (write_en==1'b1)
			r_32_31 <= data_in;
	if (addr_selector[32]&addr_selector[32])
		data_out <= r_32_32;
		if (write_en==1'b1)
			r_32_32 <= data_in;
	if (addr_selector[32]&addr_selector[33])
		data_out <= r_32_33;
		if (write_en==1'b1)
			r_32_33 <= data_in;
	if (addr_selector[32]&addr_selector[34])
		data_out <= r_32_34;
		if (write_en==1'b1)
			r_32_34 <= data_in;
	if (addr_selector[32]&addr_selector[35])
		data_out <= r_32_35;
		if (write_en==1'b1)
			r_32_35 <= data_in;
	if (addr_selector[32]&addr_selector[36])
		data_out <= r_32_36;
		if (write_en==1'b1)
			r_32_36 <= data_in;
	if (addr_selector[32]&addr_selector[37])
		data_out <= r_32_37;
		if (write_en==1'b1)
			r_32_37 <= data_in;
	if (addr_selector[32]&addr_selector[38])
		data_out <= r_32_38;
		if (write_en==1'b1)
			r_32_38 <= data_in;
	if (addr_selector[32]&addr_selector[39])
		data_out <= r_32_39;
		if (write_en==1'b1)
			r_32_39 <= data_in;
	if (addr_selector[32]&addr_selector[40])
		data_out <= r_32_40;
		if (write_en==1'b1)
			r_32_40 <= data_in;
	if (addr_selector[32]&addr_selector[41])
		data_out <= r_32_41;
		if (write_en==1'b1)
			r_32_41 <= data_in;
	if (addr_selector[32]&addr_selector[42])
		data_out <= r_32_42;
		if (write_en==1'b1)
			r_32_42 <= data_in;
	if (addr_selector[32]&addr_selector[43])
		data_out <= r_32_43;
		if (write_en==1'b1)
			r_32_43 <= data_in;
	if (addr_selector[32]&addr_selector[44])
		data_out <= r_32_44;
		if (write_en==1'b1)
			r_32_44 <= data_in;
	if (addr_selector[32]&addr_selector[45])
		data_out <= r_32_45;
		if (write_en==1'b1)
			r_32_45 <= data_in;
	if (addr_selector[32]&addr_selector[46])
		data_out <= r_32_46;
		if (write_en==1'b1)
			r_32_46 <= data_in;
	if (addr_selector[32]&addr_selector[47])
		data_out <= r_32_47;
		if (write_en==1'b1)
			r_32_47 <= data_in;
	if (addr_selector[32]&addr_selector[48])
		data_out <= r_32_48;
		if (write_en==1'b1)
			r_32_48 <= data_in;
	if (addr_selector[32]&addr_selector[49])
		data_out <= r_32_49;
		if (write_en==1'b1)
			r_32_49 <= data_in;
	if (addr_selector[32]&addr_selector[50])
		data_out <= r_32_50;
		if (write_en==1'b1)
			r_32_50 <= data_in;
	if (addr_selector[32]&addr_selector[51])
		data_out <= r_32_51;
		if (write_en==1'b1)
			r_32_51 <= data_in;
	if (addr_selector[32]&addr_selector[52])
		data_out <= r_32_52;
		if (write_en==1'b1)
			r_32_52 <= data_in;
	if (addr_selector[32]&addr_selector[53])
		data_out <= r_32_53;
		if (write_en==1'b1)
			r_32_53 <= data_in;
	if (addr_selector[32]&addr_selector[54])
		data_out <= r_32_54;
		if (write_en==1'b1)
			r_32_54 <= data_in;
	if (addr_selector[32]&addr_selector[55])
		data_out <= r_32_55;
		if (write_en==1'b1)
			r_32_55 <= data_in;
	if (addr_selector[32]&addr_selector[56])
		data_out <= r_32_56;
		if (write_en==1'b1)
			r_32_56 <= data_in;
	if (addr_selector[32]&addr_selector[57])
		data_out <= r_32_57;
		if (write_en==1'b1)
			r_32_57 <= data_in;
	if (addr_selector[32]&addr_selector[58])
		data_out <= r_32_58;
		if (write_en==1'b1)
			r_32_58 <= data_in;
	if (addr_selector[32]&addr_selector[59])
		data_out <= r_32_59;
		if (write_en==1'b1)
			r_32_59 <= data_in;
	if (addr_selector[32]&addr_selector[60])
		data_out <= r_32_60;
		if (write_en==1'b1)
			r_32_60 <= data_in;
	if (addr_selector[32]&addr_selector[61])
		data_out <= r_32_61;
		if (write_en==1'b1)
			r_32_61 <= data_in;
	if (addr_selector[32]&addr_selector[62])
		data_out <= r_32_62;
		if (write_en==1'b1)
			r_32_62 <= data_in;
	if (addr_selector[32]&addr_selector[63])
		data_out <= r_32_63;
		if (write_en==1'b1)
			r_32_63 <= data_in;
	if (addr_selector[33]&addr_selector[0])
		data_out <= r_33_0;
		if (write_en==1'b1)
			r_33_0 <= data_in;
	if (addr_selector[33]&addr_selector[1])
		data_out <= r_33_1;
		if (write_en==1'b1)
			r_33_1 <= data_in;
	if (addr_selector[33]&addr_selector[2])
		data_out <= r_33_2;
		if (write_en==1'b1)
			r_33_2 <= data_in;
	if (addr_selector[33]&addr_selector[3])
		data_out <= r_33_3;
		if (write_en==1'b1)
			r_33_3 <= data_in;
	if (addr_selector[33]&addr_selector[4])
		data_out <= r_33_4;
		if (write_en==1'b1)
			r_33_4 <= data_in;
	if (addr_selector[33]&addr_selector[5])
		data_out <= r_33_5;
		if (write_en==1'b1)
			r_33_5 <= data_in;
	if (addr_selector[33]&addr_selector[6])
		data_out <= r_33_6;
		if (write_en==1'b1)
			r_33_6 <= data_in;
	if (addr_selector[33]&addr_selector[7])
		data_out <= r_33_7;
		if (write_en==1'b1)
			r_33_7 <= data_in;
	if (addr_selector[33]&addr_selector[8])
		data_out <= r_33_8;
		if (write_en==1'b1)
			r_33_8 <= data_in;
	if (addr_selector[33]&addr_selector[9])
		data_out <= r_33_9;
		if (write_en==1'b1)
			r_33_9 <= data_in;
	if (addr_selector[33]&addr_selector[10])
		data_out <= r_33_10;
		if (write_en==1'b1)
			r_33_10 <= data_in;
	if (addr_selector[33]&addr_selector[11])
		data_out <= r_33_11;
		if (write_en==1'b1)
			r_33_11 <= data_in;
	if (addr_selector[33]&addr_selector[12])
		data_out <= r_33_12;
		if (write_en==1'b1)
			r_33_12 <= data_in;
	if (addr_selector[33]&addr_selector[13])
		data_out <= r_33_13;
		if (write_en==1'b1)
			r_33_13 <= data_in;
	if (addr_selector[33]&addr_selector[14])
		data_out <= r_33_14;
		if (write_en==1'b1)
			r_33_14 <= data_in;
	if (addr_selector[33]&addr_selector[15])
		data_out <= r_33_15;
		if (write_en==1'b1)
			r_33_15 <= data_in;
	if (addr_selector[33]&addr_selector[16])
		data_out <= r_33_16;
		if (write_en==1'b1)
			r_33_16 <= data_in;
	if (addr_selector[33]&addr_selector[17])
		data_out <= r_33_17;
		if (write_en==1'b1)
			r_33_17 <= data_in;
	if (addr_selector[33]&addr_selector[18])
		data_out <= r_33_18;
		if (write_en==1'b1)
			r_33_18 <= data_in;
	if (addr_selector[33]&addr_selector[19])
		data_out <= r_33_19;
		if (write_en==1'b1)
			r_33_19 <= data_in;
	if (addr_selector[33]&addr_selector[20])
		data_out <= r_33_20;
		if (write_en==1'b1)
			r_33_20 <= data_in;
	if (addr_selector[33]&addr_selector[21])
		data_out <= r_33_21;
		if (write_en==1'b1)
			r_33_21 <= data_in;
	if (addr_selector[33]&addr_selector[22])
		data_out <= r_33_22;
		if (write_en==1'b1)
			r_33_22 <= data_in;
	if (addr_selector[33]&addr_selector[23])
		data_out <= r_33_23;
		if (write_en==1'b1)
			r_33_23 <= data_in;
	if (addr_selector[33]&addr_selector[24])
		data_out <= r_33_24;
		if (write_en==1'b1)
			r_33_24 <= data_in;
	if (addr_selector[33]&addr_selector[25])
		data_out <= r_33_25;
		if (write_en==1'b1)
			r_33_25 <= data_in;
	if (addr_selector[33]&addr_selector[26])
		data_out <= r_33_26;
		if (write_en==1'b1)
			r_33_26 <= data_in;
	if (addr_selector[33]&addr_selector[27])
		data_out <= r_33_27;
		if (write_en==1'b1)
			r_33_27 <= data_in;
	if (addr_selector[33]&addr_selector[28])
		data_out <= r_33_28;
		if (write_en==1'b1)
			r_33_28 <= data_in;
	if (addr_selector[33]&addr_selector[29])
		data_out <= r_33_29;
		if (write_en==1'b1)
			r_33_29 <= data_in;
	if (addr_selector[33]&addr_selector[30])
		data_out <= r_33_30;
		if (write_en==1'b1)
			r_33_30 <= data_in;
	if (addr_selector[33]&addr_selector[31])
		data_out <= r_33_31;
		if (write_en==1'b1)
			r_33_31 <= data_in;
	if (addr_selector[33]&addr_selector[32])
		data_out <= r_33_32;
		if (write_en==1'b1)
			r_33_32 <= data_in;
	if (addr_selector[33]&addr_selector[33])
		data_out <= r_33_33;
		if (write_en==1'b1)
			r_33_33 <= data_in;
	if (addr_selector[33]&addr_selector[34])
		data_out <= r_33_34;
		if (write_en==1'b1)
			r_33_34 <= data_in;
	if (addr_selector[33]&addr_selector[35])
		data_out <= r_33_35;
		if (write_en==1'b1)
			r_33_35 <= data_in;
	if (addr_selector[33]&addr_selector[36])
		data_out <= r_33_36;
		if (write_en==1'b1)
			r_33_36 <= data_in;
	if (addr_selector[33]&addr_selector[37])
		data_out <= r_33_37;
		if (write_en==1'b1)
			r_33_37 <= data_in;
	if (addr_selector[33]&addr_selector[38])
		data_out <= r_33_38;
		if (write_en==1'b1)
			r_33_38 <= data_in;
	if (addr_selector[33]&addr_selector[39])
		data_out <= r_33_39;
		if (write_en==1'b1)
			r_33_39 <= data_in;
	if (addr_selector[33]&addr_selector[40])
		data_out <= r_33_40;
		if (write_en==1'b1)
			r_33_40 <= data_in;
	if (addr_selector[33]&addr_selector[41])
		data_out <= r_33_41;
		if (write_en==1'b1)
			r_33_41 <= data_in;
	if (addr_selector[33]&addr_selector[42])
		data_out <= r_33_42;
		if (write_en==1'b1)
			r_33_42 <= data_in;
	if (addr_selector[33]&addr_selector[43])
		data_out <= r_33_43;
		if (write_en==1'b1)
			r_33_43 <= data_in;
	if (addr_selector[33]&addr_selector[44])
		data_out <= r_33_44;
		if (write_en==1'b1)
			r_33_44 <= data_in;
	if (addr_selector[33]&addr_selector[45])
		data_out <= r_33_45;
		if (write_en==1'b1)
			r_33_45 <= data_in;
	if (addr_selector[33]&addr_selector[46])
		data_out <= r_33_46;
		if (write_en==1'b1)
			r_33_46 <= data_in;
	if (addr_selector[33]&addr_selector[47])
		data_out <= r_33_47;
		if (write_en==1'b1)
			r_33_47 <= data_in;
	if (addr_selector[33]&addr_selector[48])
		data_out <= r_33_48;
		if (write_en==1'b1)
			r_33_48 <= data_in;
	if (addr_selector[33]&addr_selector[49])
		data_out <= r_33_49;
		if (write_en==1'b1)
			r_33_49 <= data_in;
	if (addr_selector[33]&addr_selector[50])
		data_out <= r_33_50;
		if (write_en==1'b1)
			r_33_50 <= data_in;
	if (addr_selector[33]&addr_selector[51])
		data_out <= r_33_51;
		if (write_en==1'b1)
			r_33_51 <= data_in;
	if (addr_selector[33]&addr_selector[52])
		data_out <= r_33_52;
		if (write_en==1'b1)
			r_33_52 <= data_in;
	if (addr_selector[33]&addr_selector[53])
		data_out <= r_33_53;
		if (write_en==1'b1)
			r_33_53 <= data_in;
	if (addr_selector[33]&addr_selector[54])
		data_out <= r_33_54;
		if (write_en==1'b1)
			r_33_54 <= data_in;
	if (addr_selector[33]&addr_selector[55])
		data_out <= r_33_55;
		if (write_en==1'b1)
			r_33_55 <= data_in;
	if (addr_selector[33]&addr_selector[56])
		data_out <= r_33_56;
		if (write_en==1'b1)
			r_33_56 <= data_in;
	if (addr_selector[33]&addr_selector[57])
		data_out <= r_33_57;
		if (write_en==1'b1)
			r_33_57 <= data_in;
	if (addr_selector[33]&addr_selector[58])
		data_out <= r_33_58;
		if (write_en==1'b1)
			r_33_58 <= data_in;
	if (addr_selector[33]&addr_selector[59])
		data_out <= r_33_59;
		if (write_en==1'b1)
			r_33_59 <= data_in;
	if (addr_selector[33]&addr_selector[60])
		data_out <= r_33_60;
		if (write_en==1'b1)
			r_33_60 <= data_in;
	if (addr_selector[33]&addr_selector[61])
		data_out <= r_33_61;
		if (write_en==1'b1)
			r_33_61 <= data_in;
	if (addr_selector[33]&addr_selector[62])
		data_out <= r_33_62;
		if (write_en==1'b1)
			r_33_62 <= data_in;
	if (addr_selector[33]&addr_selector[63])
		data_out <= r_33_63;
		if (write_en==1'b1)
			r_33_63 <= data_in;
	if (addr_selector[34]&addr_selector[0])
		data_out <= r_34_0;
		if (write_en==1'b1)
			r_34_0 <= data_in;
	if (addr_selector[34]&addr_selector[1])
		data_out <= r_34_1;
		if (write_en==1'b1)
			r_34_1 <= data_in;
	if (addr_selector[34]&addr_selector[2])
		data_out <= r_34_2;
		if (write_en==1'b1)
			r_34_2 <= data_in;
	if (addr_selector[34]&addr_selector[3])
		data_out <= r_34_3;
		if (write_en==1'b1)
			r_34_3 <= data_in;
	if (addr_selector[34]&addr_selector[4])
		data_out <= r_34_4;
		if (write_en==1'b1)
			r_34_4 <= data_in;
	if (addr_selector[34]&addr_selector[5])
		data_out <= r_34_5;
		if (write_en==1'b1)
			r_34_5 <= data_in;
	if (addr_selector[34]&addr_selector[6])
		data_out <= r_34_6;
		if (write_en==1'b1)
			r_34_6 <= data_in;
	if (addr_selector[34]&addr_selector[7])
		data_out <= r_34_7;
		if (write_en==1'b1)
			r_34_7 <= data_in;
	if (addr_selector[34]&addr_selector[8])
		data_out <= r_34_8;
		if (write_en==1'b1)
			r_34_8 <= data_in;
	if (addr_selector[34]&addr_selector[9])
		data_out <= r_34_9;
		if (write_en==1'b1)
			r_34_9 <= data_in;
	if (addr_selector[34]&addr_selector[10])
		data_out <= r_34_10;
		if (write_en==1'b1)
			r_34_10 <= data_in;
	if (addr_selector[34]&addr_selector[11])
		data_out <= r_34_11;
		if (write_en==1'b1)
			r_34_11 <= data_in;
	if (addr_selector[34]&addr_selector[12])
		data_out <= r_34_12;
		if (write_en==1'b1)
			r_34_12 <= data_in;
	if (addr_selector[34]&addr_selector[13])
		data_out <= r_34_13;
		if (write_en==1'b1)
			r_34_13 <= data_in;
	if (addr_selector[34]&addr_selector[14])
		data_out <= r_34_14;
		if (write_en==1'b1)
			r_34_14 <= data_in;
	if (addr_selector[34]&addr_selector[15])
		data_out <= r_34_15;
		if (write_en==1'b1)
			r_34_15 <= data_in;
	if (addr_selector[34]&addr_selector[16])
		data_out <= r_34_16;
		if (write_en==1'b1)
			r_34_16 <= data_in;
	if (addr_selector[34]&addr_selector[17])
		data_out <= r_34_17;
		if (write_en==1'b1)
			r_34_17 <= data_in;
	if (addr_selector[34]&addr_selector[18])
		data_out <= r_34_18;
		if (write_en==1'b1)
			r_34_18 <= data_in;
	if (addr_selector[34]&addr_selector[19])
		data_out <= r_34_19;
		if (write_en==1'b1)
			r_34_19 <= data_in;
	if (addr_selector[34]&addr_selector[20])
		data_out <= r_34_20;
		if (write_en==1'b1)
			r_34_20 <= data_in;
	if (addr_selector[34]&addr_selector[21])
		data_out <= r_34_21;
		if (write_en==1'b1)
			r_34_21 <= data_in;
	if (addr_selector[34]&addr_selector[22])
		data_out <= r_34_22;
		if (write_en==1'b1)
			r_34_22 <= data_in;
	if (addr_selector[34]&addr_selector[23])
		data_out <= r_34_23;
		if (write_en==1'b1)
			r_34_23 <= data_in;
	if (addr_selector[34]&addr_selector[24])
		data_out <= r_34_24;
		if (write_en==1'b1)
			r_34_24 <= data_in;
	if (addr_selector[34]&addr_selector[25])
		data_out <= r_34_25;
		if (write_en==1'b1)
			r_34_25 <= data_in;
	if (addr_selector[34]&addr_selector[26])
		data_out <= r_34_26;
		if (write_en==1'b1)
			r_34_26 <= data_in;
	if (addr_selector[34]&addr_selector[27])
		data_out <= r_34_27;
		if (write_en==1'b1)
			r_34_27 <= data_in;
	if (addr_selector[34]&addr_selector[28])
		data_out <= r_34_28;
		if (write_en==1'b1)
			r_34_28 <= data_in;
	if (addr_selector[34]&addr_selector[29])
		data_out <= r_34_29;
		if (write_en==1'b1)
			r_34_29 <= data_in;
	if (addr_selector[34]&addr_selector[30])
		data_out <= r_34_30;
		if (write_en==1'b1)
			r_34_30 <= data_in;
	if (addr_selector[34]&addr_selector[31])
		data_out <= r_34_31;
		if (write_en==1'b1)
			r_34_31 <= data_in;
	if (addr_selector[34]&addr_selector[32])
		data_out <= r_34_32;
		if (write_en==1'b1)
			r_34_32 <= data_in;
	if (addr_selector[34]&addr_selector[33])
		data_out <= r_34_33;
		if (write_en==1'b1)
			r_34_33 <= data_in;
	if (addr_selector[34]&addr_selector[34])
		data_out <= r_34_34;
		if (write_en==1'b1)
			r_34_34 <= data_in;
	if (addr_selector[34]&addr_selector[35])
		data_out <= r_34_35;
		if (write_en==1'b1)
			r_34_35 <= data_in;
	if (addr_selector[34]&addr_selector[36])
		data_out <= r_34_36;
		if (write_en==1'b1)
			r_34_36 <= data_in;
	if (addr_selector[34]&addr_selector[37])
		data_out <= r_34_37;
		if (write_en==1'b1)
			r_34_37 <= data_in;
	if (addr_selector[34]&addr_selector[38])
		data_out <= r_34_38;
		if (write_en==1'b1)
			r_34_38 <= data_in;
	if (addr_selector[34]&addr_selector[39])
		data_out <= r_34_39;
		if (write_en==1'b1)
			r_34_39 <= data_in;
	if (addr_selector[34]&addr_selector[40])
		data_out <= r_34_40;
		if (write_en==1'b1)
			r_34_40 <= data_in;
	if (addr_selector[34]&addr_selector[41])
		data_out <= r_34_41;
		if (write_en==1'b1)
			r_34_41 <= data_in;
	if (addr_selector[34]&addr_selector[42])
		data_out <= r_34_42;
		if (write_en==1'b1)
			r_34_42 <= data_in;
	if (addr_selector[34]&addr_selector[43])
		data_out <= r_34_43;
		if (write_en==1'b1)
			r_34_43 <= data_in;
	if (addr_selector[34]&addr_selector[44])
		data_out <= r_34_44;
		if (write_en==1'b1)
			r_34_44 <= data_in;
	if (addr_selector[34]&addr_selector[45])
		data_out <= r_34_45;
		if (write_en==1'b1)
			r_34_45 <= data_in;
	if (addr_selector[34]&addr_selector[46])
		data_out <= r_34_46;
		if (write_en==1'b1)
			r_34_46 <= data_in;
	if (addr_selector[34]&addr_selector[47])
		data_out <= r_34_47;
		if (write_en==1'b1)
			r_34_47 <= data_in;
	if (addr_selector[34]&addr_selector[48])
		data_out <= r_34_48;
		if (write_en==1'b1)
			r_34_48 <= data_in;
	if (addr_selector[34]&addr_selector[49])
		data_out <= r_34_49;
		if (write_en==1'b1)
			r_34_49 <= data_in;
	if (addr_selector[34]&addr_selector[50])
		data_out <= r_34_50;
		if (write_en==1'b1)
			r_34_50 <= data_in;
	if (addr_selector[34]&addr_selector[51])
		data_out <= r_34_51;
		if (write_en==1'b1)
			r_34_51 <= data_in;
	if (addr_selector[34]&addr_selector[52])
		data_out <= r_34_52;
		if (write_en==1'b1)
			r_34_52 <= data_in;
	if (addr_selector[34]&addr_selector[53])
		data_out <= r_34_53;
		if (write_en==1'b1)
			r_34_53 <= data_in;
	if (addr_selector[34]&addr_selector[54])
		data_out <= r_34_54;
		if (write_en==1'b1)
			r_34_54 <= data_in;
	if (addr_selector[34]&addr_selector[55])
		data_out <= r_34_55;
		if (write_en==1'b1)
			r_34_55 <= data_in;
	if (addr_selector[34]&addr_selector[56])
		data_out <= r_34_56;
		if (write_en==1'b1)
			r_34_56 <= data_in;
	if (addr_selector[34]&addr_selector[57])
		data_out <= r_34_57;
		if (write_en==1'b1)
			r_34_57 <= data_in;
	if (addr_selector[34]&addr_selector[58])
		data_out <= r_34_58;
		if (write_en==1'b1)
			r_34_58 <= data_in;
	if (addr_selector[34]&addr_selector[59])
		data_out <= r_34_59;
		if (write_en==1'b1)
			r_34_59 <= data_in;
	if (addr_selector[34]&addr_selector[60])
		data_out <= r_34_60;
		if (write_en==1'b1)
			r_34_60 <= data_in;
	if (addr_selector[34]&addr_selector[61])
		data_out <= r_34_61;
		if (write_en==1'b1)
			r_34_61 <= data_in;
	if (addr_selector[34]&addr_selector[62])
		data_out <= r_34_62;
		if (write_en==1'b1)
			r_34_62 <= data_in;
	if (addr_selector[34]&addr_selector[63])
		data_out <= r_34_63;
		if (write_en==1'b1)
			r_34_63 <= data_in;
	if (addr_selector[35]&addr_selector[0])
		data_out <= r_35_0;
		if (write_en==1'b1)
			r_35_0 <= data_in;
	if (addr_selector[35]&addr_selector[1])
		data_out <= r_35_1;
		if (write_en==1'b1)
			r_35_1 <= data_in;
	if (addr_selector[35]&addr_selector[2])
		data_out <= r_35_2;
		if (write_en==1'b1)
			r_35_2 <= data_in;
	if (addr_selector[35]&addr_selector[3])
		data_out <= r_35_3;
		if (write_en==1'b1)
			r_35_3 <= data_in;
	if (addr_selector[35]&addr_selector[4])
		data_out <= r_35_4;
		if (write_en==1'b1)
			r_35_4 <= data_in;
	if (addr_selector[35]&addr_selector[5])
		data_out <= r_35_5;
		if (write_en==1'b1)
			r_35_5 <= data_in;
	if (addr_selector[35]&addr_selector[6])
		data_out <= r_35_6;
		if (write_en==1'b1)
			r_35_6 <= data_in;
	if (addr_selector[35]&addr_selector[7])
		data_out <= r_35_7;
		if (write_en==1'b1)
			r_35_7 <= data_in;
	if (addr_selector[35]&addr_selector[8])
		data_out <= r_35_8;
		if (write_en==1'b1)
			r_35_8 <= data_in;
	if (addr_selector[35]&addr_selector[9])
		data_out <= r_35_9;
		if (write_en==1'b1)
			r_35_9 <= data_in;
	if (addr_selector[35]&addr_selector[10])
		data_out <= r_35_10;
		if (write_en==1'b1)
			r_35_10 <= data_in;
	if (addr_selector[35]&addr_selector[11])
		data_out <= r_35_11;
		if (write_en==1'b1)
			r_35_11 <= data_in;
	if (addr_selector[35]&addr_selector[12])
		data_out <= r_35_12;
		if (write_en==1'b1)
			r_35_12 <= data_in;
	if (addr_selector[35]&addr_selector[13])
		data_out <= r_35_13;
		if (write_en==1'b1)
			r_35_13 <= data_in;
	if (addr_selector[35]&addr_selector[14])
		data_out <= r_35_14;
		if (write_en==1'b1)
			r_35_14 <= data_in;
	if (addr_selector[35]&addr_selector[15])
		data_out <= r_35_15;
		if (write_en==1'b1)
			r_35_15 <= data_in;
	if (addr_selector[35]&addr_selector[16])
		data_out <= r_35_16;
		if (write_en==1'b1)
			r_35_16 <= data_in;
	if (addr_selector[35]&addr_selector[17])
		data_out <= r_35_17;
		if (write_en==1'b1)
			r_35_17 <= data_in;
	if (addr_selector[35]&addr_selector[18])
		data_out <= r_35_18;
		if (write_en==1'b1)
			r_35_18 <= data_in;
	if (addr_selector[35]&addr_selector[19])
		data_out <= r_35_19;
		if (write_en==1'b1)
			r_35_19 <= data_in;
	if (addr_selector[35]&addr_selector[20])
		data_out <= r_35_20;
		if (write_en==1'b1)
			r_35_20 <= data_in;
	if (addr_selector[35]&addr_selector[21])
		data_out <= r_35_21;
		if (write_en==1'b1)
			r_35_21 <= data_in;
	if (addr_selector[35]&addr_selector[22])
		data_out <= r_35_22;
		if (write_en==1'b1)
			r_35_22 <= data_in;
	if (addr_selector[35]&addr_selector[23])
		data_out <= r_35_23;
		if (write_en==1'b1)
			r_35_23 <= data_in;
	if (addr_selector[35]&addr_selector[24])
		data_out <= r_35_24;
		if (write_en==1'b1)
			r_35_24 <= data_in;
	if (addr_selector[35]&addr_selector[25])
		data_out <= r_35_25;
		if (write_en==1'b1)
			r_35_25 <= data_in;
	if (addr_selector[35]&addr_selector[26])
		data_out <= r_35_26;
		if (write_en==1'b1)
			r_35_26 <= data_in;
	if (addr_selector[35]&addr_selector[27])
		data_out <= r_35_27;
		if (write_en==1'b1)
			r_35_27 <= data_in;
	if (addr_selector[35]&addr_selector[28])
		data_out <= r_35_28;
		if (write_en==1'b1)
			r_35_28 <= data_in;
	if (addr_selector[35]&addr_selector[29])
		data_out <= r_35_29;
		if (write_en==1'b1)
			r_35_29 <= data_in;
	if (addr_selector[35]&addr_selector[30])
		data_out <= r_35_30;
		if (write_en==1'b1)
			r_35_30 <= data_in;
	if (addr_selector[35]&addr_selector[31])
		data_out <= r_35_31;
		if (write_en==1'b1)
			r_35_31 <= data_in;
	if (addr_selector[35]&addr_selector[32])
		data_out <= r_35_32;
		if (write_en==1'b1)
			r_35_32 <= data_in;
	if (addr_selector[35]&addr_selector[33])
		data_out <= r_35_33;
		if (write_en==1'b1)
			r_35_33 <= data_in;
	if (addr_selector[35]&addr_selector[34])
		data_out <= r_35_34;
		if (write_en==1'b1)
			r_35_34 <= data_in;
	if (addr_selector[35]&addr_selector[35])
		data_out <= r_35_35;
		if (write_en==1'b1)
			r_35_35 <= data_in;
	if (addr_selector[35]&addr_selector[36])
		data_out <= r_35_36;
		if (write_en==1'b1)
			r_35_36 <= data_in;
	if (addr_selector[35]&addr_selector[37])
		data_out <= r_35_37;
		if (write_en==1'b1)
			r_35_37 <= data_in;
	if (addr_selector[35]&addr_selector[38])
		data_out <= r_35_38;
		if (write_en==1'b1)
			r_35_38 <= data_in;
	if (addr_selector[35]&addr_selector[39])
		data_out <= r_35_39;
		if (write_en==1'b1)
			r_35_39 <= data_in;
	if (addr_selector[35]&addr_selector[40])
		data_out <= r_35_40;
		if (write_en==1'b1)
			r_35_40 <= data_in;
	if (addr_selector[35]&addr_selector[41])
		data_out <= r_35_41;
		if (write_en==1'b1)
			r_35_41 <= data_in;
	if (addr_selector[35]&addr_selector[42])
		data_out <= r_35_42;
		if (write_en==1'b1)
			r_35_42 <= data_in;
	if (addr_selector[35]&addr_selector[43])
		data_out <= r_35_43;
		if (write_en==1'b1)
			r_35_43 <= data_in;
	if (addr_selector[35]&addr_selector[44])
		data_out <= r_35_44;
		if (write_en==1'b1)
			r_35_44 <= data_in;
	if (addr_selector[35]&addr_selector[45])
		data_out <= r_35_45;
		if (write_en==1'b1)
			r_35_45 <= data_in;
	if (addr_selector[35]&addr_selector[46])
		data_out <= r_35_46;
		if (write_en==1'b1)
			r_35_46 <= data_in;
	if (addr_selector[35]&addr_selector[47])
		data_out <= r_35_47;
		if (write_en==1'b1)
			r_35_47 <= data_in;
	if (addr_selector[35]&addr_selector[48])
		data_out <= r_35_48;
		if (write_en==1'b1)
			r_35_48 <= data_in;
	if (addr_selector[35]&addr_selector[49])
		data_out <= r_35_49;
		if (write_en==1'b1)
			r_35_49 <= data_in;
	if (addr_selector[35]&addr_selector[50])
		data_out <= r_35_50;
		if (write_en==1'b1)
			r_35_50 <= data_in;
	if (addr_selector[35]&addr_selector[51])
		data_out <= r_35_51;
		if (write_en==1'b1)
			r_35_51 <= data_in;
	if (addr_selector[35]&addr_selector[52])
		data_out <= r_35_52;
		if (write_en==1'b1)
			r_35_52 <= data_in;
	if (addr_selector[35]&addr_selector[53])
		data_out <= r_35_53;
		if (write_en==1'b1)
			r_35_53 <= data_in;
	if (addr_selector[35]&addr_selector[54])
		data_out <= r_35_54;
		if (write_en==1'b1)
			r_35_54 <= data_in;
	if (addr_selector[35]&addr_selector[55])
		data_out <= r_35_55;
		if (write_en==1'b1)
			r_35_55 <= data_in;
	if (addr_selector[35]&addr_selector[56])
		data_out <= r_35_56;
		if (write_en==1'b1)
			r_35_56 <= data_in;
	if (addr_selector[35]&addr_selector[57])
		data_out <= r_35_57;
		if (write_en==1'b1)
			r_35_57 <= data_in;
	if (addr_selector[35]&addr_selector[58])
		data_out <= r_35_58;
		if (write_en==1'b1)
			r_35_58 <= data_in;
	if (addr_selector[35]&addr_selector[59])
		data_out <= r_35_59;
		if (write_en==1'b1)
			r_35_59 <= data_in;
	if (addr_selector[35]&addr_selector[60])
		data_out <= r_35_60;
		if (write_en==1'b1)
			r_35_60 <= data_in;
	if (addr_selector[35]&addr_selector[61])
		data_out <= r_35_61;
		if (write_en==1'b1)
			r_35_61 <= data_in;
	if (addr_selector[35]&addr_selector[62])
		data_out <= r_35_62;
		if (write_en==1'b1)
			r_35_62 <= data_in;
	if (addr_selector[35]&addr_selector[63])
		data_out <= r_35_63;
		if (write_en==1'b1)
			r_35_63 <= data_in;
	if (addr_selector[36]&addr_selector[0])
		data_out <= r_36_0;
		if (write_en==1'b1)
			r_36_0 <= data_in;
	if (addr_selector[36]&addr_selector[1])
		data_out <= r_36_1;
		if (write_en==1'b1)
			r_36_1 <= data_in;
	if (addr_selector[36]&addr_selector[2])
		data_out <= r_36_2;
		if (write_en==1'b1)
			r_36_2 <= data_in;
	if (addr_selector[36]&addr_selector[3])
		data_out <= r_36_3;
		if (write_en==1'b1)
			r_36_3 <= data_in;
	if (addr_selector[36]&addr_selector[4])
		data_out <= r_36_4;
		if (write_en==1'b1)
			r_36_4 <= data_in;
	if (addr_selector[36]&addr_selector[5])
		data_out <= r_36_5;
		if (write_en==1'b1)
			r_36_5 <= data_in;
	if (addr_selector[36]&addr_selector[6])
		data_out <= r_36_6;
		if (write_en==1'b1)
			r_36_6 <= data_in;
	if (addr_selector[36]&addr_selector[7])
		data_out <= r_36_7;
		if (write_en==1'b1)
			r_36_7 <= data_in;
	if (addr_selector[36]&addr_selector[8])
		data_out <= r_36_8;
		if (write_en==1'b1)
			r_36_8 <= data_in;
	if (addr_selector[36]&addr_selector[9])
		data_out <= r_36_9;
		if (write_en==1'b1)
			r_36_9 <= data_in;
	if (addr_selector[36]&addr_selector[10])
		data_out <= r_36_10;
		if (write_en==1'b1)
			r_36_10 <= data_in;
	if (addr_selector[36]&addr_selector[11])
		data_out <= r_36_11;
		if (write_en==1'b1)
			r_36_11 <= data_in;
	if (addr_selector[36]&addr_selector[12])
		data_out <= r_36_12;
		if (write_en==1'b1)
			r_36_12 <= data_in;
	if (addr_selector[36]&addr_selector[13])
		data_out <= r_36_13;
		if (write_en==1'b1)
			r_36_13 <= data_in;
	if (addr_selector[36]&addr_selector[14])
		data_out <= r_36_14;
		if (write_en==1'b1)
			r_36_14 <= data_in;
	if (addr_selector[36]&addr_selector[15])
		data_out <= r_36_15;
		if (write_en==1'b1)
			r_36_15 <= data_in;
	if (addr_selector[36]&addr_selector[16])
		data_out <= r_36_16;
		if (write_en==1'b1)
			r_36_16 <= data_in;
	if (addr_selector[36]&addr_selector[17])
		data_out <= r_36_17;
		if (write_en==1'b1)
			r_36_17 <= data_in;
	if (addr_selector[36]&addr_selector[18])
		data_out <= r_36_18;
		if (write_en==1'b1)
			r_36_18 <= data_in;
	if (addr_selector[36]&addr_selector[19])
		data_out <= r_36_19;
		if (write_en==1'b1)
			r_36_19 <= data_in;
	if (addr_selector[36]&addr_selector[20])
		data_out <= r_36_20;
		if (write_en==1'b1)
			r_36_20 <= data_in;
	if (addr_selector[36]&addr_selector[21])
		data_out <= r_36_21;
		if (write_en==1'b1)
			r_36_21 <= data_in;
	if (addr_selector[36]&addr_selector[22])
		data_out <= r_36_22;
		if (write_en==1'b1)
			r_36_22 <= data_in;
	if (addr_selector[36]&addr_selector[23])
		data_out <= r_36_23;
		if (write_en==1'b1)
			r_36_23 <= data_in;
	if (addr_selector[36]&addr_selector[24])
		data_out <= r_36_24;
		if (write_en==1'b1)
			r_36_24 <= data_in;
	if (addr_selector[36]&addr_selector[25])
		data_out <= r_36_25;
		if (write_en==1'b1)
			r_36_25 <= data_in;
	if (addr_selector[36]&addr_selector[26])
		data_out <= r_36_26;
		if (write_en==1'b1)
			r_36_26 <= data_in;
	if (addr_selector[36]&addr_selector[27])
		data_out <= r_36_27;
		if (write_en==1'b1)
			r_36_27 <= data_in;
	if (addr_selector[36]&addr_selector[28])
		data_out <= r_36_28;
		if (write_en==1'b1)
			r_36_28 <= data_in;
	if (addr_selector[36]&addr_selector[29])
		data_out <= r_36_29;
		if (write_en==1'b1)
			r_36_29 <= data_in;
	if (addr_selector[36]&addr_selector[30])
		data_out <= r_36_30;
		if (write_en==1'b1)
			r_36_30 <= data_in;
	if (addr_selector[36]&addr_selector[31])
		data_out <= r_36_31;
		if (write_en==1'b1)
			r_36_31 <= data_in;
	if (addr_selector[36]&addr_selector[32])
		data_out <= r_36_32;
		if (write_en==1'b1)
			r_36_32 <= data_in;
	if (addr_selector[36]&addr_selector[33])
		data_out <= r_36_33;
		if (write_en==1'b1)
			r_36_33 <= data_in;
	if (addr_selector[36]&addr_selector[34])
		data_out <= r_36_34;
		if (write_en==1'b1)
			r_36_34 <= data_in;
	if (addr_selector[36]&addr_selector[35])
		data_out <= r_36_35;
		if (write_en==1'b1)
			r_36_35 <= data_in;
	if (addr_selector[36]&addr_selector[36])
		data_out <= r_36_36;
		if (write_en==1'b1)
			r_36_36 <= data_in;
	if (addr_selector[36]&addr_selector[37])
		data_out <= r_36_37;
		if (write_en==1'b1)
			r_36_37 <= data_in;
	if (addr_selector[36]&addr_selector[38])
		data_out <= r_36_38;
		if (write_en==1'b1)
			r_36_38 <= data_in;
	if (addr_selector[36]&addr_selector[39])
		data_out <= r_36_39;
		if (write_en==1'b1)
			r_36_39 <= data_in;
	if (addr_selector[36]&addr_selector[40])
		data_out <= r_36_40;
		if (write_en==1'b1)
			r_36_40 <= data_in;
	if (addr_selector[36]&addr_selector[41])
		data_out <= r_36_41;
		if (write_en==1'b1)
			r_36_41 <= data_in;
	if (addr_selector[36]&addr_selector[42])
		data_out <= r_36_42;
		if (write_en==1'b1)
			r_36_42 <= data_in;
	if (addr_selector[36]&addr_selector[43])
		data_out <= r_36_43;
		if (write_en==1'b1)
			r_36_43 <= data_in;
	if (addr_selector[36]&addr_selector[44])
		data_out <= r_36_44;
		if (write_en==1'b1)
			r_36_44 <= data_in;
	if (addr_selector[36]&addr_selector[45])
		data_out <= r_36_45;
		if (write_en==1'b1)
			r_36_45 <= data_in;
	if (addr_selector[36]&addr_selector[46])
		data_out <= r_36_46;
		if (write_en==1'b1)
			r_36_46 <= data_in;
	if (addr_selector[36]&addr_selector[47])
		data_out <= r_36_47;
		if (write_en==1'b1)
			r_36_47 <= data_in;
	if (addr_selector[36]&addr_selector[48])
		data_out <= r_36_48;
		if (write_en==1'b1)
			r_36_48 <= data_in;
	if (addr_selector[36]&addr_selector[49])
		data_out <= r_36_49;
		if (write_en==1'b1)
			r_36_49 <= data_in;
	if (addr_selector[36]&addr_selector[50])
		data_out <= r_36_50;
		if (write_en==1'b1)
			r_36_50 <= data_in;
	if (addr_selector[36]&addr_selector[51])
		data_out <= r_36_51;
		if (write_en==1'b1)
			r_36_51 <= data_in;
	if (addr_selector[36]&addr_selector[52])
		data_out <= r_36_52;
		if (write_en==1'b1)
			r_36_52 <= data_in;
	if (addr_selector[36]&addr_selector[53])
		data_out <= r_36_53;
		if (write_en==1'b1)
			r_36_53 <= data_in;
	if (addr_selector[36]&addr_selector[54])
		data_out <= r_36_54;
		if (write_en==1'b1)
			r_36_54 <= data_in;
	if (addr_selector[36]&addr_selector[55])
		data_out <= r_36_55;
		if (write_en==1'b1)
			r_36_55 <= data_in;
	if (addr_selector[36]&addr_selector[56])
		data_out <= r_36_56;
		if (write_en==1'b1)
			r_36_56 <= data_in;
	if (addr_selector[36]&addr_selector[57])
		data_out <= r_36_57;
		if (write_en==1'b1)
			r_36_57 <= data_in;
	if (addr_selector[36]&addr_selector[58])
		data_out <= r_36_58;
		if (write_en==1'b1)
			r_36_58 <= data_in;
	if (addr_selector[36]&addr_selector[59])
		data_out <= r_36_59;
		if (write_en==1'b1)
			r_36_59 <= data_in;
	if (addr_selector[36]&addr_selector[60])
		data_out <= r_36_60;
		if (write_en==1'b1)
			r_36_60 <= data_in;
	if (addr_selector[36]&addr_selector[61])
		data_out <= r_36_61;
		if (write_en==1'b1)
			r_36_61 <= data_in;
	if (addr_selector[36]&addr_selector[62])
		data_out <= r_36_62;
		if (write_en==1'b1)
			r_36_62 <= data_in;
	if (addr_selector[36]&addr_selector[63])
		data_out <= r_36_63;
		if (write_en==1'b1)
			r_36_63 <= data_in;
	if (addr_selector[37]&addr_selector[0])
		data_out <= r_37_0;
		if (write_en==1'b1)
			r_37_0 <= data_in;
	if (addr_selector[37]&addr_selector[1])
		data_out <= r_37_1;
		if (write_en==1'b1)
			r_37_1 <= data_in;
	if (addr_selector[37]&addr_selector[2])
		data_out <= r_37_2;
		if (write_en==1'b1)
			r_37_2 <= data_in;
	if (addr_selector[37]&addr_selector[3])
		data_out <= r_37_3;
		if (write_en==1'b1)
			r_37_3 <= data_in;
	if (addr_selector[37]&addr_selector[4])
		data_out <= r_37_4;
		if (write_en==1'b1)
			r_37_4 <= data_in;
	if (addr_selector[37]&addr_selector[5])
		data_out <= r_37_5;
		if (write_en==1'b1)
			r_37_5 <= data_in;
	if (addr_selector[37]&addr_selector[6])
		data_out <= r_37_6;
		if (write_en==1'b1)
			r_37_6 <= data_in;
	if (addr_selector[37]&addr_selector[7])
		data_out <= r_37_7;
		if (write_en==1'b1)
			r_37_7 <= data_in;
	if (addr_selector[37]&addr_selector[8])
		data_out <= r_37_8;
		if (write_en==1'b1)
			r_37_8 <= data_in;
	if (addr_selector[37]&addr_selector[9])
		data_out <= r_37_9;
		if (write_en==1'b1)
			r_37_9 <= data_in;
	if (addr_selector[37]&addr_selector[10])
		data_out <= r_37_10;
		if (write_en==1'b1)
			r_37_10 <= data_in;
	if (addr_selector[37]&addr_selector[11])
		data_out <= r_37_11;
		if (write_en==1'b1)
			r_37_11 <= data_in;
	if (addr_selector[37]&addr_selector[12])
		data_out <= r_37_12;
		if (write_en==1'b1)
			r_37_12 <= data_in;
	if (addr_selector[37]&addr_selector[13])
		data_out <= r_37_13;
		if (write_en==1'b1)
			r_37_13 <= data_in;
	if (addr_selector[37]&addr_selector[14])
		data_out <= r_37_14;
		if (write_en==1'b1)
			r_37_14 <= data_in;
	if (addr_selector[37]&addr_selector[15])
		data_out <= r_37_15;
		if (write_en==1'b1)
			r_37_15 <= data_in;
	if (addr_selector[37]&addr_selector[16])
		data_out <= r_37_16;
		if (write_en==1'b1)
			r_37_16 <= data_in;
	if (addr_selector[37]&addr_selector[17])
		data_out <= r_37_17;
		if (write_en==1'b1)
			r_37_17 <= data_in;
	if (addr_selector[37]&addr_selector[18])
		data_out <= r_37_18;
		if (write_en==1'b1)
			r_37_18 <= data_in;
	if (addr_selector[37]&addr_selector[19])
		data_out <= r_37_19;
		if (write_en==1'b1)
			r_37_19 <= data_in;
	if (addr_selector[37]&addr_selector[20])
		data_out <= r_37_20;
		if (write_en==1'b1)
			r_37_20 <= data_in;
	if (addr_selector[37]&addr_selector[21])
		data_out <= r_37_21;
		if (write_en==1'b1)
			r_37_21 <= data_in;
	if (addr_selector[37]&addr_selector[22])
		data_out <= r_37_22;
		if (write_en==1'b1)
			r_37_22 <= data_in;
	if (addr_selector[37]&addr_selector[23])
		data_out <= r_37_23;
		if (write_en==1'b1)
			r_37_23 <= data_in;
	if (addr_selector[37]&addr_selector[24])
		data_out <= r_37_24;
		if (write_en==1'b1)
			r_37_24 <= data_in;
	if (addr_selector[37]&addr_selector[25])
		data_out <= r_37_25;
		if (write_en==1'b1)
			r_37_25 <= data_in;
	if (addr_selector[37]&addr_selector[26])
		data_out <= r_37_26;
		if (write_en==1'b1)
			r_37_26 <= data_in;
	if (addr_selector[37]&addr_selector[27])
		data_out <= r_37_27;
		if (write_en==1'b1)
			r_37_27 <= data_in;
	if (addr_selector[37]&addr_selector[28])
		data_out <= r_37_28;
		if (write_en==1'b1)
			r_37_28 <= data_in;
	if (addr_selector[37]&addr_selector[29])
		data_out <= r_37_29;
		if (write_en==1'b1)
			r_37_29 <= data_in;
	if (addr_selector[37]&addr_selector[30])
		data_out <= r_37_30;
		if (write_en==1'b1)
			r_37_30 <= data_in;
	if (addr_selector[37]&addr_selector[31])
		data_out <= r_37_31;
		if (write_en==1'b1)
			r_37_31 <= data_in;
	if (addr_selector[37]&addr_selector[32])
		data_out <= r_37_32;
		if (write_en==1'b1)
			r_37_32 <= data_in;
	if (addr_selector[37]&addr_selector[33])
		data_out <= r_37_33;
		if (write_en==1'b1)
			r_37_33 <= data_in;
	if (addr_selector[37]&addr_selector[34])
		data_out <= r_37_34;
		if (write_en==1'b1)
			r_37_34 <= data_in;
	if (addr_selector[37]&addr_selector[35])
		data_out <= r_37_35;
		if (write_en==1'b1)
			r_37_35 <= data_in;
	if (addr_selector[37]&addr_selector[36])
		data_out <= r_37_36;
		if (write_en==1'b1)
			r_37_36 <= data_in;
	if (addr_selector[37]&addr_selector[37])
		data_out <= r_37_37;
		if (write_en==1'b1)
			r_37_37 <= data_in;
	if (addr_selector[37]&addr_selector[38])
		data_out <= r_37_38;
		if (write_en==1'b1)
			r_37_38 <= data_in;
	if (addr_selector[37]&addr_selector[39])
		data_out <= r_37_39;
		if (write_en==1'b1)
			r_37_39 <= data_in;
	if (addr_selector[37]&addr_selector[40])
		data_out <= r_37_40;
		if (write_en==1'b1)
			r_37_40 <= data_in;
	if (addr_selector[37]&addr_selector[41])
		data_out <= r_37_41;
		if (write_en==1'b1)
			r_37_41 <= data_in;
	if (addr_selector[37]&addr_selector[42])
		data_out <= r_37_42;
		if (write_en==1'b1)
			r_37_42 <= data_in;
	if (addr_selector[37]&addr_selector[43])
		data_out <= r_37_43;
		if (write_en==1'b1)
			r_37_43 <= data_in;
	if (addr_selector[37]&addr_selector[44])
		data_out <= r_37_44;
		if (write_en==1'b1)
			r_37_44 <= data_in;
	if (addr_selector[37]&addr_selector[45])
		data_out <= r_37_45;
		if (write_en==1'b1)
			r_37_45 <= data_in;
	if (addr_selector[37]&addr_selector[46])
		data_out <= r_37_46;
		if (write_en==1'b1)
			r_37_46 <= data_in;
	if (addr_selector[37]&addr_selector[47])
		data_out <= r_37_47;
		if (write_en==1'b1)
			r_37_47 <= data_in;
	if (addr_selector[37]&addr_selector[48])
		data_out <= r_37_48;
		if (write_en==1'b1)
			r_37_48 <= data_in;
	if (addr_selector[37]&addr_selector[49])
		data_out <= r_37_49;
		if (write_en==1'b1)
			r_37_49 <= data_in;
	if (addr_selector[37]&addr_selector[50])
		data_out <= r_37_50;
		if (write_en==1'b1)
			r_37_50 <= data_in;
	if (addr_selector[37]&addr_selector[51])
		data_out <= r_37_51;
		if (write_en==1'b1)
			r_37_51 <= data_in;
	if (addr_selector[37]&addr_selector[52])
		data_out <= r_37_52;
		if (write_en==1'b1)
			r_37_52 <= data_in;
	if (addr_selector[37]&addr_selector[53])
		data_out <= r_37_53;
		if (write_en==1'b1)
			r_37_53 <= data_in;
	if (addr_selector[37]&addr_selector[54])
		data_out <= r_37_54;
		if (write_en==1'b1)
			r_37_54 <= data_in;
	if (addr_selector[37]&addr_selector[55])
		data_out <= r_37_55;
		if (write_en==1'b1)
			r_37_55 <= data_in;
	if (addr_selector[37]&addr_selector[56])
		data_out <= r_37_56;
		if (write_en==1'b1)
			r_37_56 <= data_in;
	if (addr_selector[37]&addr_selector[57])
		data_out <= r_37_57;
		if (write_en==1'b1)
			r_37_57 <= data_in;
	if (addr_selector[37]&addr_selector[58])
		data_out <= r_37_58;
		if (write_en==1'b1)
			r_37_58 <= data_in;
	if (addr_selector[37]&addr_selector[59])
		data_out <= r_37_59;
		if (write_en==1'b1)
			r_37_59 <= data_in;
	if (addr_selector[37]&addr_selector[60])
		data_out <= r_37_60;
		if (write_en==1'b1)
			r_37_60 <= data_in;
	if (addr_selector[37]&addr_selector[61])
		data_out <= r_37_61;
		if (write_en==1'b1)
			r_37_61 <= data_in;
	if (addr_selector[37]&addr_selector[62])
		data_out <= r_37_62;
		if (write_en==1'b1)
			r_37_62 <= data_in;
	if (addr_selector[37]&addr_selector[63])
		data_out <= r_37_63;
		if (write_en==1'b1)
			r_37_63 <= data_in;
	if (addr_selector[38]&addr_selector[0])
		data_out <= r_38_0;
		if (write_en==1'b1)
			r_38_0 <= data_in;
	if (addr_selector[38]&addr_selector[1])
		data_out <= r_38_1;
		if (write_en==1'b1)
			r_38_1 <= data_in;
	if (addr_selector[38]&addr_selector[2])
		data_out <= r_38_2;
		if (write_en==1'b1)
			r_38_2 <= data_in;
	if (addr_selector[38]&addr_selector[3])
		data_out <= r_38_3;
		if (write_en==1'b1)
			r_38_3 <= data_in;
	if (addr_selector[38]&addr_selector[4])
		data_out <= r_38_4;
		if (write_en==1'b1)
			r_38_4 <= data_in;
	if (addr_selector[38]&addr_selector[5])
		data_out <= r_38_5;
		if (write_en==1'b1)
			r_38_5 <= data_in;
	if (addr_selector[38]&addr_selector[6])
		data_out <= r_38_6;
		if (write_en==1'b1)
			r_38_6 <= data_in;
	if (addr_selector[38]&addr_selector[7])
		data_out <= r_38_7;
		if (write_en==1'b1)
			r_38_7 <= data_in;
	if (addr_selector[38]&addr_selector[8])
		data_out <= r_38_8;
		if (write_en==1'b1)
			r_38_8 <= data_in;
	if (addr_selector[38]&addr_selector[9])
		data_out <= r_38_9;
		if (write_en==1'b1)
			r_38_9 <= data_in;
	if (addr_selector[38]&addr_selector[10])
		data_out <= r_38_10;
		if (write_en==1'b1)
			r_38_10 <= data_in;
	if (addr_selector[38]&addr_selector[11])
		data_out <= r_38_11;
		if (write_en==1'b1)
			r_38_11 <= data_in;
	if (addr_selector[38]&addr_selector[12])
		data_out <= r_38_12;
		if (write_en==1'b1)
			r_38_12 <= data_in;
	if (addr_selector[38]&addr_selector[13])
		data_out <= r_38_13;
		if (write_en==1'b1)
			r_38_13 <= data_in;
	if (addr_selector[38]&addr_selector[14])
		data_out <= r_38_14;
		if (write_en==1'b1)
			r_38_14 <= data_in;
	if (addr_selector[38]&addr_selector[15])
		data_out <= r_38_15;
		if (write_en==1'b1)
			r_38_15 <= data_in;
	if (addr_selector[38]&addr_selector[16])
		data_out <= r_38_16;
		if (write_en==1'b1)
			r_38_16 <= data_in;
	if (addr_selector[38]&addr_selector[17])
		data_out <= r_38_17;
		if (write_en==1'b1)
			r_38_17 <= data_in;
	if (addr_selector[38]&addr_selector[18])
		data_out <= r_38_18;
		if (write_en==1'b1)
			r_38_18 <= data_in;
	if (addr_selector[38]&addr_selector[19])
		data_out <= r_38_19;
		if (write_en==1'b1)
			r_38_19 <= data_in;
	if (addr_selector[38]&addr_selector[20])
		data_out <= r_38_20;
		if (write_en==1'b1)
			r_38_20 <= data_in;
	if (addr_selector[38]&addr_selector[21])
		data_out <= r_38_21;
		if (write_en==1'b1)
			r_38_21 <= data_in;
	if (addr_selector[38]&addr_selector[22])
		data_out <= r_38_22;
		if (write_en==1'b1)
			r_38_22 <= data_in;
	if (addr_selector[38]&addr_selector[23])
		data_out <= r_38_23;
		if (write_en==1'b1)
			r_38_23 <= data_in;
	if (addr_selector[38]&addr_selector[24])
		data_out <= r_38_24;
		if (write_en==1'b1)
			r_38_24 <= data_in;
	if (addr_selector[38]&addr_selector[25])
		data_out <= r_38_25;
		if (write_en==1'b1)
			r_38_25 <= data_in;
	if (addr_selector[38]&addr_selector[26])
		data_out <= r_38_26;
		if (write_en==1'b1)
			r_38_26 <= data_in;
	if (addr_selector[38]&addr_selector[27])
		data_out <= r_38_27;
		if (write_en==1'b1)
			r_38_27 <= data_in;
	if (addr_selector[38]&addr_selector[28])
		data_out <= r_38_28;
		if (write_en==1'b1)
			r_38_28 <= data_in;
	if (addr_selector[38]&addr_selector[29])
		data_out <= r_38_29;
		if (write_en==1'b1)
			r_38_29 <= data_in;
	if (addr_selector[38]&addr_selector[30])
		data_out <= r_38_30;
		if (write_en==1'b1)
			r_38_30 <= data_in;
	if (addr_selector[38]&addr_selector[31])
		data_out <= r_38_31;
		if (write_en==1'b1)
			r_38_31 <= data_in;
	if (addr_selector[38]&addr_selector[32])
		data_out <= r_38_32;
		if (write_en==1'b1)
			r_38_32 <= data_in;
	if (addr_selector[38]&addr_selector[33])
		data_out <= r_38_33;
		if (write_en==1'b1)
			r_38_33 <= data_in;
	if (addr_selector[38]&addr_selector[34])
		data_out <= r_38_34;
		if (write_en==1'b1)
			r_38_34 <= data_in;
	if (addr_selector[38]&addr_selector[35])
		data_out <= r_38_35;
		if (write_en==1'b1)
			r_38_35 <= data_in;
	if (addr_selector[38]&addr_selector[36])
		data_out <= r_38_36;
		if (write_en==1'b1)
			r_38_36 <= data_in;
	if (addr_selector[38]&addr_selector[37])
		data_out <= r_38_37;
		if (write_en==1'b1)
			r_38_37 <= data_in;
	if (addr_selector[38]&addr_selector[38])
		data_out <= r_38_38;
		if (write_en==1'b1)
			r_38_38 <= data_in;
	if (addr_selector[38]&addr_selector[39])
		data_out <= r_38_39;
		if (write_en==1'b1)
			r_38_39 <= data_in;
	if (addr_selector[38]&addr_selector[40])
		data_out <= r_38_40;
		if (write_en==1'b1)
			r_38_40 <= data_in;
	if (addr_selector[38]&addr_selector[41])
		data_out <= r_38_41;
		if (write_en==1'b1)
			r_38_41 <= data_in;
	if (addr_selector[38]&addr_selector[42])
		data_out <= r_38_42;
		if (write_en==1'b1)
			r_38_42 <= data_in;
	if (addr_selector[38]&addr_selector[43])
		data_out <= r_38_43;
		if (write_en==1'b1)
			r_38_43 <= data_in;
	if (addr_selector[38]&addr_selector[44])
		data_out <= r_38_44;
		if (write_en==1'b1)
			r_38_44 <= data_in;
	if (addr_selector[38]&addr_selector[45])
		data_out <= r_38_45;
		if (write_en==1'b1)
			r_38_45 <= data_in;
	if (addr_selector[38]&addr_selector[46])
		data_out <= r_38_46;
		if (write_en==1'b1)
			r_38_46 <= data_in;
	if (addr_selector[38]&addr_selector[47])
		data_out <= r_38_47;
		if (write_en==1'b1)
			r_38_47 <= data_in;
	if (addr_selector[38]&addr_selector[48])
		data_out <= r_38_48;
		if (write_en==1'b1)
			r_38_48 <= data_in;
	if (addr_selector[38]&addr_selector[49])
		data_out <= r_38_49;
		if (write_en==1'b1)
			r_38_49 <= data_in;
	if (addr_selector[38]&addr_selector[50])
		data_out <= r_38_50;
		if (write_en==1'b1)
			r_38_50 <= data_in;
	if (addr_selector[38]&addr_selector[51])
		data_out <= r_38_51;
		if (write_en==1'b1)
			r_38_51 <= data_in;
	if (addr_selector[38]&addr_selector[52])
		data_out <= r_38_52;
		if (write_en==1'b1)
			r_38_52 <= data_in;
	if (addr_selector[38]&addr_selector[53])
		data_out <= r_38_53;
		if (write_en==1'b1)
			r_38_53 <= data_in;
	if (addr_selector[38]&addr_selector[54])
		data_out <= r_38_54;
		if (write_en==1'b1)
			r_38_54 <= data_in;
	if (addr_selector[38]&addr_selector[55])
		data_out <= r_38_55;
		if (write_en==1'b1)
			r_38_55 <= data_in;
	if (addr_selector[38]&addr_selector[56])
		data_out <= r_38_56;
		if (write_en==1'b1)
			r_38_56 <= data_in;
	if (addr_selector[38]&addr_selector[57])
		data_out <= r_38_57;
		if (write_en==1'b1)
			r_38_57 <= data_in;
	if (addr_selector[38]&addr_selector[58])
		data_out <= r_38_58;
		if (write_en==1'b1)
			r_38_58 <= data_in;
	if (addr_selector[38]&addr_selector[59])
		data_out <= r_38_59;
		if (write_en==1'b1)
			r_38_59 <= data_in;
	if (addr_selector[38]&addr_selector[60])
		data_out <= r_38_60;
		if (write_en==1'b1)
			r_38_60 <= data_in;
	if (addr_selector[38]&addr_selector[61])
		data_out <= r_38_61;
		if (write_en==1'b1)
			r_38_61 <= data_in;
	if (addr_selector[38]&addr_selector[62])
		data_out <= r_38_62;
		if (write_en==1'b1)
			r_38_62 <= data_in;
	if (addr_selector[38]&addr_selector[63])
		data_out <= r_38_63;
		if (write_en==1'b1)
			r_38_63 <= data_in;
	if (addr_selector[39]&addr_selector[0])
		data_out <= r_39_0;
		if (write_en==1'b1)
			r_39_0 <= data_in;
	if (addr_selector[39]&addr_selector[1])
		data_out <= r_39_1;
		if (write_en==1'b1)
			r_39_1 <= data_in;
	if (addr_selector[39]&addr_selector[2])
		data_out <= r_39_2;
		if (write_en==1'b1)
			r_39_2 <= data_in;
	if (addr_selector[39]&addr_selector[3])
		data_out <= r_39_3;
		if (write_en==1'b1)
			r_39_3 <= data_in;
	if (addr_selector[39]&addr_selector[4])
		data_out <= r_39_4;
		if (write_en==1'b1)
			r_39_4 <= data_in;
	if (addr_selector[39]&addr_selector[5])
		data_out <= r_39_5;
		if (write_en==1'b1)
			r_39_5 <= data_in;
	if (addr_selector[39]&addr_selector[6])
		data_out <= r_39_6;
		if (write_en==1'b1)
			r_39_6 <= data_in;
	if (addr_selector[39]&addr_selector[7])
		data_out <= r_39_7;
		if (write_en==1'b1)
			r_39_7 <= data_in;
	if (addr_selector[39]&addr_selector[8])
		data_out <= r_39_8;
		if (write_en==1'b1)
			r_39_8 <= data_in;
	if (addr_selector[39]&addr_selector[9])
		data_out <= r_39_9;
		if (write_en==1'b1)
			r_39_9 <= data_in;
	if (addr_selector[39]&addr_selector[10])
		data_out <= r_39_10;
		if (write_en==1'b1)
			r_39_10 <= data_in;
	if (addr_selector[39]&addr_selector[11])
		data_out <= r_39_11;
		if (write_en==1'b1)
			r_39_11 <= data_in;
	if (addr_selector[39]&addr_selector[12])
		data_out <= r_39_12;
		if (write_en==1'b1)
			r_39_12 <= data_in;
	if (addr_selector[39]&addr_selector[13])
		data_out <= r_39_13;
		if (write_en==1'b1)
			r_39_13 <= data_in;
	if (addr_selector[39]&addr_selector[14])
		data_out <= r_39_14;
		if (write_en==1'b1)
			r_39_14 <= data_in;
	if (addr_selector[39]&addr_selector[15])
		data_out <= r_39_15;
		if (write_en==1'b1)
			r_39_15 <= data_in;
	if (addr_selector[39]&addr_selector[16])
		data_out <= r_39_16;
		if (write_en==1'b1)
			r_39_16 <= data_in;
	if (addr_selector[39]&addr_selector[17])
		data_out <= r_39_17;
		if (write_en==1'b1)
			r_39_17 <= data_in;
	if (addr_selector[39]&addr_selector[18])
		data_out <= r_39_18;
		if (write_en==1'b1)
			r_39_18 <= data_in;
	if (addr_selector[39]&addr_selector[19])
		data_out <= r_39_19;
		if (write_en==1'b1)
			r_39_19 <= data_in;
	if (addr_selector[39]&addr_selector[20])
		data_out <= r_39_20;
		if (write_en==1'b1)
			r_39_20 <= data_in;
	if (addr_selector[39]&addr_selector[21])
		data_out <= r_39_21;
		if (write_en==1'b1)
			r_39_21 <= data_in;
	if (addr_selector[39]&addr_selector[22])
		data_out <= r_39_22;
		if (write_en==1'b1)
			r_39_22 <= data_in;
	if (addr_selector[39]&addr_selector[23])
		data_out <= r_39_23;
		if (write_en==1'b1)
			r_39_23 <= data_in;
	if (addr_selector[39]&addr_selector[24])
		data_out <= r_39_24;
		if (write_en==1'b1)
			r_39_24 <= data_in;
	if (addr_selector[39]&addr_selector[25])
		data_out <= r_39_25;
		if (write_en==1'b1)
			r_39_25 <= data_in;
	if (addr_selector[39]&addr_selector[26])
		data_out <= r_39_26;
		if (write_en==1'b1)
			r_39_26 <= data_in;
	if (addr_selector[39]&addr_selector[27])
		data_out <= r_39_27;
		if (write_en==1'b1)
			r_39_27 <= data_in;
	if (addr_selector[39]&addr_selector[28])
		data_out <= r_39_28;
		if (write_en==1'b1)
			r_39_28 <= data_in;
	if (addr_selector[39]&addr_selector[29])
		data_out <= r_39_29;
		if (write_en==1'b1)
			r_39_29 <= data_in;
	if (addr_selector[39]&addr_selector[30])
		data_out <= r_39_30;
		if (write_en==1'b1)
			r_39_30 <= data_in;
	if (addr_selector[39]&addr_selector[31])
		data_out <= r_39_31;
		if (write_en==1'b1)
			r_39_31 <= data_in;
	if (addr_selector[39]&addr_selector[32])
		data_out <= r_39_32;
		if (write_en==1'b1)
			r_39_32 <= data_in;
	if (addr_selector[39]&addr_selector[33])
		data_out <= r_39_33;
		if (write_en==1'b1)
			r_39_33 <= data_in;
	if (addr_selector[39]&addr_selector[34])
		data_out <= r_39_34;
		if (write_en==1'b1)
			r_39_34 <= data_in;
	if (addr_selector[39]&addr_selector[35])
		data_out <= r_39_35;
		if (write_en==1'b1)
			r_39_35 <= data_in;
	if (addr_selector[39]&addr_selector[36])
		data_out <= r_39_36;
		if (write_en==1'b1)
			r_39_36 <= data_in;
	if (addr_selector[39]&addr_selector[37])
		data_out <= r_39_37;
		if (write_en==1'b1)
			r_39_37 <= data_in;
	if (addr_selector[39]&addr_selector[38])
		data_out <= r_39_38;
		if (write_en==1'b1)
			r_39_38 <= data_in;
	if (addr_selector[39]&addr_selector[39])
		data_out <= r_39_39;
		if (write_en==1'b1)
			r_39_39 <= data_in;
	if (addr_selector[39]&addr_selector[40])
		data_out <= r_39_40;
		if (write_en==1'b1)
			r_39_40 <= data_in;
	if (addr_selector[39]&addr_selector[41])
		data_out <= r_39_41;
		if (write_en==1'b1)
			r_39_41 <= data_in;
	if (addr_selector[39]&addr_selector[42])
		data_out <= r_39_42;
		if (write_en==1'b1)
			r_39_42 <= data_in;
	if (addr_selector[39]&addr_selector[43])
		data_out <= r_39_43;
		if (write_en==1'b1)
			r_39_43 <= data_in;
	if (addr_selector[39]&addr_selector[44])
		data_out <= r_39_44;
		if (write_en==1'b1)
			r_39_44 <= data_in;
	if (addr_selector[39]&addr_selector[45])
		data_out <= r_39_45;
		if (write_en==1'b1)
			r_39_45 <= data_in;
	if (addr_selector[39]&addr_selector[46])
		data_out <= r_39_46;
		if (write_en==1'b1)
			r_39_46 <= data_in;
	if (addr_selector[39]&addr_selector[47])
		data_out <= r_39_47;
		if (write_en==1'b1)
			r_39_47 <= data_in;
	if (addr_selector[39]&addr_selector[48])
		data_out <= r_39_48;
		if (write_en==1'b1)
			r_39_48 <= data_in;
	if (addr_selector[39]&addr_selector[49])
		data_out <= r_39_49;
		if (write_en==1'b1)
			r_39_49 <= data_in;
	if (addr_selector[39]&addr_selector[50])
		data_out <= r_39_50;
		if (write_en==1'b1)
			r_39_50 <= data_in;
	if (addr_selector[39]&addr_selector[51])
		data_out <= r_39_51;
		if (write_en==1'b1)
			r_39_51 <= data_in;
	if (addr_selector[39]&addr_selector[52])
		data_out <= r_39_52;
		if (write_en==1'b1)
			r_39_52 <= data_in;
	if (addr_selector[39]&addr_selector[53])
		data_out <= r_39_53;
		if (write_en==1'b1)
			r_39_53 <= data_in;
	if (addr_selector[39]&addr_selector[54])
		data_out <= r_39_54;
		if (write_en==1'b1)
			r_39_54 <= data_in;
	if (addr_selector[39]&addr_selector[55])
		data_out <= r_39_55;
		if (write_en==1'b1)
			r_39_55 <= data_in;
	if (addr_selector[39]&addr_selector[56])
		data_out <= r_39_56;
		if (write_en==1'b1)
			r_39_56 <= data_in;
	if (addr_selector[39]&addr_selector[57])
		data_out <= r_39_57;
		if (write_en==1'b1)
			r_39_57 <= data_in;
	if (addr_selector[39]&addr_selector[58])
		data_out <= r_39_58;
		if (write_en==1'b1)
			r_39_58 <= data_in;
	if (addr_selector[39]&addr_selector[59])
		data_out <= r_39_59;
		if (write_en==1'b1)
			r_39_59 <= data_in;
	if (addr_selector[39]&addr_selector[60])
		data_out <= r_39_60;
		if (write_en==1'b1)
			r_39_60 <= data_in;
	if (addr_selector[39]&addr_selector[61])
		data_out <= r_39_61;
		if (write_en==1'b1)
			r_39_61 <= data_in;
	if (addr_selector[39]&addr_selector[62])
		data_out <= r_39_62;
		if (write_en==1'b1)
			r_39_62 <= data_in;
	if (addr_selector[39]&addr_selector[63])
		data_out <= r_39_63;
		if (write_en==1'b1)
			r_39_63 <= data_in;
	if (addr_selector[40]&addr_selector[0])
		data_out <= r_40_0;
		if (write_en==1'b1)
			r_40_0 <= data_in;
	if (addr_selector[40]&addr_selector[1])
		data_out <= r_40_1;
		if (write_en==1'b1)
			r_40_1 <= data_in;
	if (addr_selector[40]&addr_selector[2])
		data_out <= r_40_2;
		if (write_en==1'b1)
			r_40_2 <= data_in;
	if (addr_selector[40]&addr_selector[3])
		data_out <= r_40_3;
		if (write_en==1'b1)
			r_40_3 <= data_in;
	if (addr_selector[40]&addr_selector[4])
		data_out <= r_40_4;
		if (write_en==1'b1)
			r_40_4 <= data_in;
	if (addr_selector[40]&addr_selector[5])
		data_out <= r_40_5;
		if (write_en==1'b1)
			r_40_5 <= data_in;
	if (addr_selector[40]&addr_selector[6])
		data_out <= r_40_6;
		if (write_en==1'b1)
			r_40_6 <= data_in;
	if (addr_selector[40]&addr_selector[7])
		data_out <= r_40_7;
		if (write_en==1'b1)
			r_40_7 <= data_in;
	if (addr_selector[40]&addr_selector[8])
		data_out <= r_40_8;
		if (write_en==1'b1)
			r_40_8 <= data_in;
	if (addr_selector[40]&addr_selector[9])
		data_out <= r_40_9;
		if (write_en==1'b1)
			r_40_9 <= data_in;
	if (addr_selector[40]&addr_selector[10])
		data_out <= r_40_10;
		if (write_en==1'b1)
			r_40_10 <= data_in;
	if (addr_selector[40]&addr_selector[11])
		data_out <= r_40_11;
		if (write_en==1'b1)
			r_40_11 <= data_in;
	if (addr_selector[40]&addr_selector[12])
		data_out <= r_40_12;
		if (write_en==1'b1)
			r_40_12 <= data_in;
	if (addr_selector[40]&addr_selector[13])
		data_out <= r_40_13;
		if (write_en==1'b1)
			r_40_13 <= data_in;
	if (addr_selector[40]&addr_selector[14])
		data_out <= r_40_14;
		if (write_en==1'b1)
			r_40_14 <= data_in;
	if (addr_selector[40]&addr_selector[15])
		data_out <= r_40_15;
		if (write_en==1'b1)
			r_40_15 <= data_in;
	if (addr_selector[40]&addr_selector[16])
		data_out <= r_40_16;
		if (write_en==1'b1)
			r_40_16 <= data_in;
	if (addr_selector[40]&addr_selector[17])
		data_out <= r_40_17;
		if (write_en==1'b1)
			r_40_17 <= data_in;
	if (addr_selector[40]&addr_selector[18])
		data_out <= r_40_18;
		if (write_en==1'b1)
			r_40_18 <= data_in;
	if (addr_selector[40]&addr_selector[19])
		data_out <= r_40_19;
		if (write_en==1'b1)
			r_40_19 <= data_in;
	if (addr_selector[40]&addr_selector[20])
		data_out <= r_40_20;
		if (write_en==1'b1)
			r_40_20 <= data_in;
	if (addr_selector[40]&addr_selector[21])
		data_out <= r_40_21;
		if (write_en==1'b1)
			r_40_21 <= data_in;
	if (addr_selector[40]&addr_selector[22])
		data_out <= r_40_22;
		if (write_en==1'b1)
			r_40_22 <= data_in;
	if (addr_selector[40]&addr_selector[23])
		data_out <= r_40_23;
		if (write_en==1'b1)
			r_40_23 <= data_in;
	if (addr_selector[40]&addr_selector[24])
		data_out <= r_40_24;
		if (write_en==1'b1)
			r_40_24 <= data_in;
	if (addr_selector[40]&addr_selector[25])
		data_out <= r_40_25;
		if (write_en==1'b1)
			r_40_25 <= data_in;
	if (addr_selector[40]&addr_selector[26])
		data_out <= r_40_26;
		if (write_en==1'b1)
			r_40_26 <= data_in;
	if (addr_selector[40]&addr_selector[27])
		data_out <= r_40_27;
		if (write_en==1'b1)
			r_40_27 <= data_in;
	if (addr_selector[40]&addr_selector[28])
		data_out <= r_40_28;
		if (write_en==1'b1)
			r_40_28 <= data_in;
	if (addr_selector[40]&addr_selector[29])
		data_out <= r_40_29;
		if (write_en==1'b1)
			r_40_29 <= data_in;
	if (addr_selector[40]&addr_selector[30])
		data_out <= r_40_30;
		if (write_en==1'b1)
			r_40_30 <= data_in;
	if (addr_selector[40]&addr_selector[31])
		data_out <= r_40_31;
		if (write_en==1'b1)
			r_40_31 <= data_in;
	if (addr_selector[40]&addr_selector[32])
		data_out <= r_40_32;
		if (write_en==1'b1)
			r_40_32 <= data_in;
	if (addr_selector[40]&addr_selector[33])
		data_out <= r_40_33;
		if (write_en==1'b1)
			r_40_33 <= data_in;
	if (addr_selector[40]&addr_selector[34])
		data_out <= r_40_34;
		if (write_en==1'b1)
			r_40_34 <= data_in;
	if (addr_selector[40]&addr_selector[35])
		data_out <= r_40_35;
		if (write_en==1'b1)
			r_40_35 <= data_in;
	if (addr_selector[40]&addr_selector[36])
		data_out <= r_40_36;
		if (write_en==1'b1)
			r_40_36 <= data_in;
	if (addr_selector[40]&addr_selector[37])
		data_out <= r_40_37;
		if (write_en==1'b1)
			r_40_37 <= data_in;
	if (addr_selector[40]&addr_selector[38])
		data_out <= r_40_38;
		if (write_en==1'b1)
			r_40_38 <= data_in;
	if (addr_selector[40]&addr_selector[39])
		data_out <= r_40_39;
		if (write_en==1'b1)
			r_40_39 <= data_in;
	if (addr_selector[40]&addr_selector[40])
		data_out <= r_40_40;
		if (write_en==1'b1)
			r_40_40 <= data_in;
	if (addr_selector[40]&addr_selector[41])
		data_out <= r_40_41;
		if (write_en==1'b1)
			r_40_41 <= data_in;
	if (addr_selector[40]&addr_selector[42])
		data_out <= r_40_42;
		if (write_en==1'b1)
			r_40_42 <= data_in;
	if (addr_selector[40]&addr_selector[43])
		data_out <= r_40_43;
		if (write_en==1'b1)
			r_40_43 <= data_in;
	if (addr_selector[40]&addr_selector[44])
		data_out <= r_40_44;
		if (write_en==1'b1)
			r_40_44 <= data_in;
	if (addr_selector[40]&addr_selector[45])
		data_out <= r_40_45;
		if (write_en==1'b1)
			r_40_45 <= data_in;
	if (addr_selector[40]&addr_selector[46])
		data_out <= r_40_46;
		if (write_en==1'b1)
			r_40_46 <= data_in;
	if (addr_selector[40]&addr_selector[47])
		data_out <= r_40_47;
		if (write_en==1'b1)
			r_40_47 <= data_in;
	if (addr_selector[40]&addr_selector[48])
		data_out <= r_40_48;
		if (write_en==1'b1)
			r_40_48 <= data_in;
	if (addr_selector[40]&addr_selector[49])
		data_out <= r_40_49;
		if (write_en==1'b1)
			r_40_49 <= data_in;
	if (addr_selector[40]&addr_selector[50])
		data_out <= r_40_50;
		if (write_en==1'b1)
			r_40_50 <= data_in;
	if (addr_selector[40]&addr_selector[51])
		data_out <= r_40_51;
		if (write_en==1'b1)
			r_40_51 <= data_in;
	if (addr_selector[40]&addr_selector[52])
		data_out <= r_40_52;
		if (write_en==1'b1)
			r_40_52 <= data_in;
	if (addr_selector[40]&addr_selector[53])
		data_out <= r_40_53;
		if (write_en==1'b1)
			r_40_53 <= data_in;
	if (addr_selector[40]&addr_selector[54])
		data_out <= r_40_54;
		if (write_en==1'b1)
			r_40_54 <= data_in;
	if (addr_selector[40]&addr_selector[55])
		data_out <= r_40_55;
		if (write_en==1'b1)
			r_40_55 <= data_in;
	if (addr_selector[40]&addr_selector[56])
		data_out <= r_40_56;
		if (write_en==1'b1)
			r_40_56 <= data_in;
	if (addr_selector[40]&addr_selector[57])
		data_out <= r_40_57;
		if (write_en==1'b1)
			r_40_57 <= data_in;
	if (addr_selector[40]&addr_selector[58])
		data_out <= r_40_58;
		if (write_en==1'b1)
			r_40_58 <= data_in;
	if (addr_selector[40]&addr_selector[59])
		data_out <= r_40_59;
		if (write_en==1'b1)
			r_40_59 <= data_in;
	if (addr_selector[40]&addr_selector[60])
		data_out <= r_40_60;
		if (write_en==1'b1)
			r_40_60 <= data_in;
	if (addr_selector[40]&addr_selector[61])
		data_out <= r_40_61;
		if (write_en==1'b1)
			r_40_61 <= data_in;
	if (addr_selector[40]&addr_selector[62])
		data_out <= r_40_62;
		if (write_en==1'b1)
			r_40_62 <= data_in;
	if (addr_selector[40]&addr_selector[63])
		data_out <= r_40_63;
		if (write_en==1'b1)
			r_40_63 <= data_in;
	if (addr_selector[41]&addr_selector[0])
		data_out <= r_41_0;
		if (write_en==1'b1)
			r_41_0 <= data_in;
	if (addr_selector[41]&addr_selector[1])
		data_out <= r_41_1;
		if (write_en==1'b1)
			r_41_1 <= data_in;
	if (addr_selector[41]&addr_selector[2])
		data_out <= r_41_2;
		if (write_en==1'b1)
			r_41_2 <= data_in;
	if (addr_selector[41]&addr_selector[3])
		data_out <= r_41_3;
		if (write_en==1'b1)
			r_41_3 <= data_in;
	if (addr_selector[41]&addr_selector[4])
		data_out <= r_41_4;
		if (write_en==1'b1)
			r_41_4 <= data_in;
	if (addr_selector[41]&addr_selector[5])
		data_out <= r_41_5;
		if (write_en==1'b1)
			r_41_5 <= data_in;
	if (addr_selector[41]&addr_selector[6])
		data_out <= r_41_6;
		if (write_en==1'b1)
			r_41_6 <= data_in;
	if (addr_selector[41]&addr_selector[7])
		data_out <= r_41_7;
		if (write_en==1'b1)
			r_41_7 <= data_in;
	if (addr_selector[41]&addr_selector[8])
		data_out <= r_41_8;
		if (write_en==1'b1)
			r_41_8 <= data_in;
	if (addr_selector[41]&addr_selector[9])
		data_out <= r_41_9;
		if (write_en==1'b1)
			r_41_9 <= data_in;
	if (addr_selector[41]&addr_selector[10])
		data_out <= r_41_10;
		if (write_en==1'b1)
			r_41_10 <= data_in;
	if (addr_selector[41]&addr_selector[11])
		data_out <= r_41_11;
		if (write_en==1'b1)
			r_41_11 <= data_in;
	if (addr_selector[41]&addr_selector[12])
		data_out <= r_41_12;
		if (write_en==1'b1)
			r_41_12 <= data_in;
	if (addr_selector[41]&addr_selector[13])
		data_out <= r_41_13;
		if (write_en==1'b1)
			r_41_13 <= data_in;
	if (addr_selector[41]&addr_selector[14])
		data_out <= r_41_14;
		if (write_en==1'b1)
			r_41_14 <= data_in;
	if (addr_selector[41]&addr_selector[15])
		data_out <= r_41_15;
		if (write_en==1'b1)
			r_41_15 <= data_in;
	if (addr_selector[41]&addr_selector[16])
		data_out <= r_41_16;
		if (write_en==1'b1)
			r_41_16 <= data_in;
	if (addr_selector[41]&addr_selector[17])
		data_out <= r_41_17;
		if (write_en==1'b1)
			r_41_17 <= data_in;
	if (addr_selector[41]&addr_selector[18])
		data_out <= r_41_18;
		if (write_en==1'b1)
			r_41_18 <= data_in;
	if (addr_selector[41]&addr_selector[19])
		data_out <= r_41_19;
		if (write_en==1'b1)
			r_41_19 <= data_in;
	if (addr_selector[41]&addr_selector[20])
		data_out <= r_41_20;
		if (write_en==1'b1)
			r_41_20 <= data_in;
	if (addr_selector[41]&addr_selector[21])
		data_out <= r_41_21;
		if (write_en==1'b1)
			r_41_21 <= data_in;
	if (addr_selector[41]&addr_selector[22])
		data_out <= r_41_22;
		if (write_en==1'b1)
			r_41_22 <= data_in;
	if (addr_selector[41]&addr_selector[23])
		data_out <= r_41_23;
		if (write_en==1'b1)
			r_41_23 <= data_in;
	if (addr_selector[41]&addr_selector[24])
		data_out <= r_41_24;
		if (write_en==1'b1)
			r_41_24 <= data_in;
	if (addr_selector[41]&addr_selector[25])
		data_out <= r_41_25;
		if (write_en==1'b1)
			r_41_25 <= data_in;
	if (addr_selector[41]&addr_selector[26])
		data_out <= r_41_26;
		if (write_en==1'b1)
			r_41_26 <= data_in;
	if (addr_selector[41]&addr_selector[27])
		data_out <= r_41_27;
		if (write_en==1'b1)
			r_41_27 <= data_in;
	if (addr_selector[41]&addr_selector[28])
		data_out <= r_41_28;
		if (write_en==1'b1)
			r_41_28 <= data_in;
	if (addr_selector[41]&addr_selector[29])
		data_out <= r_41_29;
		if (write_en==1'b1)
			r_41_29 <= data_in;
	if (addr_selector[41]&addr_selector[30])
		data_out <= r_41_30;
		if (write_en==1'b1)
			r_41_30 <= data_in;
	if (addr_selector[41]&addr_selector[31])
		data_out <= r_41_31;
		if (write_en==1'b1)
			r_41_31 <= data_in;
	if (addr_selector[41]&addr_selector[32])
		data_out <= r_41_32;
		if (write_en==1'b1)
			r_41_32 <= data_in;
	if (addr_selector[41]&addr_selector[33])
		data_out <= r_41_33;
		if (write_en==1'b1)
			r_41_33 <= data_in;
	if (addr_selector[41]&addr_selector[34])
		data_out <= r_41_34;
		if (write_en==1'b1)
			r_41_34 <= data_in;
	if (addr_selector[41]&addr_selector[35])
		data_out <= r_41_35;
		if (write_en==1'b1)
			r_41_35 <= data_in;
	if (addr_selector[41]&addr_selector[36])
		data_out <= r_41_36;
		if (write_en==1'b1)
			r_41_36 <= data_in;
	if (addr_selector[41]&addr_selector[37])
		data_out <= r_41_37;
		if (write_en==1'b1)
			r_41_37 <= data_in;
	if (addr_selector[41]&addr_selector[38])
		data_out <= r_41_38;
		if (write_en==1'b1)
			r_41_38 <= data_in;
	if (addr_selector[41]&addr_selector[39])
		data_out <= r_41_39;
		if (write_en==1'b1)
			r_41_39 <= data_in;
	if (addr_selector[41]&addr_selector[40])
		data_out <= r_41_40;
		if (write_en==1'b1)
			r_41_40 <= data_in;
	if (addr_selector[41]&addr_selector[41])
		data_out <= r_41_41;
		if (write_en==1'b1)
			r_41_41 <= data_in;
	if (addr_selector[41]&addr_selector[42])
		data_out <= r_41_42;
		if (write_en==1'b1)
			r_41_42 <= data_in;
	if (addr_selector[41]&addr_selector[43])
		data_out <= r_41_43;
		if (write_en==1'b1)
			r_41_43 <= data_in;
	if (addr_selector[41]&addr_selector[44])
		data_out <= r_41_44;
		if (write_en==1'b1)
			r_41_44 <= data_in;
	if (addr_selector[41]&addr_selector[45])
		data_out <= r_41_45;
		if (write_en==1'b1)
			r_41_45 <= data_in;
	if (addr_selector[41]&addr_selector[46])
		data_out <= r_41_46;
		if (write_en==1'b1)
			r_41_46 <= data_in;
	if (addr_selector[41]&addr_selector[47])
		data_out <= r_41_47;
		if (write_en==1'b1)
			r_41_47 <= data_in;
	if (addr_selector[41]&addr_selector[48])
		data_out <= r_41_48;
		if (write_en==1'b1)
			r_41_48 <= data_in;
	if (addr_selector[41]&addr_selector[49])
		data_out <= r_41_49;
		if (write_en==1'b1)
			r_41_49 <= data_in;
	if (addr_selector[41]&addr_selector[50])
		data_out <= r_41_50;
		if (write_en==1'b1)
			r_41_50 <= data_in;
	if (addr_selector[41]&addr_selector[51])
		data_out <= r_41_51;
		if (write_en==1'b1)
			r_41_51 <= data_in;
	if (addr_selector[41]&addr_selector[52])
		data_out <= r_41_52;
		if (write_en==1'b1)
			r_41_52 <= data_in;
	if (addr_selector[41]&addr_selector[53])
		data_out <= r_41_53;
		if (write_en==1'b1)
			r_41_53 <= data_in;
	if (addr_selector[41]&addr_selector[54])
		data_out <= r_41_54;
		if (write_en==1'b1)
			r_41_54 <= data_in;
	if (addr_selector[41]&addr_selector[55])
		data_out <= r_41_55;
		if (write_en==1'b1)
			r_41_55 <= data_in;
	if (addr_selector[41]&addr_selector[56])
		data_out <= r_41_56;
		if (write_en==1'b1)
			r_41_56 <= data_in;
	if (addr_selector[41]&addr_selector[57])
		data_out <= r_41_57;
		if (write_en==1'b1)
			r_41_57 <= data_in;
	if (addr_selector[41]&addr_selector[58])
		data_out <= r_41_58;
		if (write_en==1'b1)
			r_41_58 <= data_in;
	if (addr_selector[41]&addr_selector[59])
		data_out <= r_41_59;
		if (write_en==1'b1)
			r_41_59 <= data_in;
	if (addr_selector[41]&addr_selector[60])
		data_out <= r_41_60;
		if (write_en==1'b1)
			r_41_60 <= data_in;
	if (addr_selector[41]&addr_selector[61])
		data_out <= r_41_61;
		if (write_en==1'b1)
			r_41_61 <= data_in;
	if (addr_selector[41]&addr_selector[62])
		data_out <= r_41_62;
		if (write_en==1'b1)
			r_41_62 <= data_in;
	if (addr_selector[41]&addr_selector[63])
		data_out <= r_41_63;
		if (write_en==1'b1)
			r_41_63 <= data_in;
	if (addr_selector[42]&addr_selector[0])
		data_out <= r_42_0;
		if (write_en==1'b1)
			r_42_0 <= data_in;
	if (addr_selector[42]&addr_selector[1])
		data_out <= r_42_1;
		if (write_en==1'b1)
			r_42_1 <= data_in;
	if (addr_selector[42]&addr_selector[2])
		data_out <= r_42_2;
		if (write_en==1'b1)
			r_42_2 <= data_in;
	if (addr_selector[42]&addr_selector[3])
		data_out <= r_42_3;
		if (write_en==1'b1)
			r_42_3 <= data_in;
	if (addr_selector[42]&addr_selector[4])
		data_out <= r_42_4;
		if (write_en==1'b1)
			r_42_4 <= data_in;
	if (addr_selector[42]&addr_selector[5])
		data_out <= r_42_5;
		if (write_en==1'b1)
			r_42_5 <= data_in;
	if (addr_selector[42]&addr_selector[6])
		data_out <= r_42_6;
		if (write_en==1'b1)
			r_42_6 <= data_in;
	if (addr_selector[42]&addr_selector[7])
		data_out <= r_42_7;
		if (write_en==1'b1)
			r_42_7 <= data_in;
	if (addr_selector[42]&addr_selector[8])
		data_out <= r_42_8;
		if (write_en==1'b1)
			r_42_8 <= data_in;
	if (addr_selector[42]&addr_selector[9])
		data_out <= r_42_9;
		if (write_en==1'b1)
			r_42_9 <= data_in;
	if (addr_selector[42]&addr_selector[10])
		data_out <= r_42_10;
		if (write_en==1'b1)
			r_42_10 <= data_in;
	if (addr_selector[42]&addr_selector[11])
		data_out <= r_42_11;
		if (write_en==1'b1)
			r_42_11 <= data_in;
	if (addr_selector[42]&addr_selector[12])
		data_out <= r_42_12;
		if (write_en==1'b1)
			r_42_12 <= data_in;
	if (addr_selector[42]&addr_selector[13])
		data_out <= r_42_13;
		if (write_en==1'b1)
			r_42_13 <= data_in;
	if (addr_selector[42]&addr_selector[14])
		data_out <= r_42_14;
		if (write_en==1'b1)
			r_42_14 <= data_in;
	if (addr_selector[42]&addr_selector[15])
		data_out <= r_42_15;
		if (write_en==1'b1)
			r_42_15 <= data_in;
	if (addr_selector[42]&addr_selector[16])
		data_out <= r_42_16;
		if (write_en==1'b1)
			r_42_16 <= data_in;
	if (addr_selector[42]&addr_selector[17])
		data_out <= r_42_17;
		if (write_en==1'b1)
			r_42_17 <= data_in;
	if (addr_selector[42]&addr_selector[18])
		data_out <= r_42_18;
		if (write_en==1'b1)
			r_42_18 <= data_in;
	if (addr_selector[42]&addr_selector[19])
		data_out <= r_42_19;
		if (write_en==1'b1)
			r_42_19 <= data_in;
	if (addr_selector[42]&addr_selector[20])
		data_out <= r_42_20;
		if (write_en==1'b1)
			r_42_20 <= data_in;
	if (addr_selector[42]&addr_selector[21])
		data_out <= r_42_21;
		if (write_en==1'b1)
			r_42_21 <= data_in;
	if (addr_selector[42]&addr_selector[22])
		data_out <= r_42_22;
		if (write_en==1'b1)
			r_42_22 <= data_in;
	if (addr_selector[42]&addr_selector[23])
		data_out <= r_42_23;
		if (write_en==1'b1)
			r_42_23 <= data_in;
	if (addr_selector[42]&addr_selector[24])
		data_out <= r_42_24;
		if (write_en==1'b1)
			r_42_24 <= data_in;
	if (addr_selector[42]&addr_selector[25])
		data_out <= r_42_25;
		if (write_en==1'b1)
			r_42_25 <= data_in;
	if (addr_selector[42]&addr_selector[26])
		data_out <= r_42_26;
		if (write_en==1'b1)
			r_42_26 <= data_in;
	if (addr_selector[42]&addr_selector[27])
		data_out <= r_42_27;
		if (write_en==1'b1)
			r_42_27 <= data_in;
	if (addr_selector[42]&addr_selector[28])
		data_out <= r_42_28;
		if (write_en==1'b1)
			r_42_28 <= data_in;
	if (addr_selector[42]&addr_selector[29])
		data_out <= r_42_29;
		if (write_en==1'b1)
			r_42_29 <= data_in;
	if (addr_selector[42]&addr_selector[30])
		data_out <= r_42_30;
		if (write_en==1'b1)
			r_42_30 <= data_in;
	if (addr_selector[42]&addr_selector[31])
		data_out <= r_42_31;
		if (write_en==1'b1)
			r_42_31 <= data_in;
	if (addr_selector[42]&addr_selector[32])
		data_out <= r_42_32;
		if (write_en==1'b1)
			r_42_32 <= data_in;
	if (addr_selector[42]&addr_selector[33])
		data_out <= r_42_33;
		if (write_en==1'b1)
			r_42_33 <= data_in;
	if (addr_selector[42]&addr_selector[34])
		data_out <= r_42_34;
		if (write_en==1'b1)
			r_42_34 <= data_in;
	if (addr_selector[42]&addr_selector[35])
		data_out <= r_42_35;
		if (write_en==1'b1)
			r_42_35 <= data_in;
	if (addr_selector[42]&addr_selector[36])
		data_out <= r_42_36;
		if (write_en==1'b1)
			r_42_36 <= data_in;
	if (addr_selector[42]&addr_selector[37])
		data_out <= r_42_37;
		if (write_en==1'b1)
			r_42_37 <= data_in;
	if (addr_selector[42]&addr_selector[38])
		data_out <= r_42_38;
		if (write_en==1'b1)
			r_42_38 <= data_in;
	if (addr_selector[42]&addr_selector[39])
		data_out <= r_42_39;
		if (write_en==1'b1)
			r_42_39 <= data_in;
	if (addr_selector[42]&addr_selector[40])
		data_out <= r_42_40;
		if (write_en==1'b1)
			r_42_40 <= data_in;
	if (addr_selector[42]&addr_selector[41])
		data_out <= r_42_41;
		if (write_en==1'b1)
			r_42_41 <= data_in;
	if (addr_selector[42]&addr_selector[42])
		data_out <= r_42_42;
		if (write_en==1'b1)
			r_42_42 <= data_in;
	if (addr_selector[42]&addr_selector[43])
		data_out <= r_42_43;
		if (write_en==1'b1)
			r_42_43 <= data_in;
	if (addr_selector[42]&addr_selector[44])
		data_out <= r_42_44;
		if (write_en==1'b1)
			r_42_44 <= data_in;
	if (addr_selector[42]&addr_selector[45])
		data_out <= r_42_45;
		if (write_en==1'b1)
			r_42_45 <= data_in;
	if (addr_selector[42]&addr_selector[46])
		data_out <= r_42_46;
		if (write_en==1'b1)
			r_42_46 <= data_in;
	if (addr_selector[42]&addr_selector[47])
		data_out <= r_42_47;
		if (write_en==1'b1)
			r_42_47 <= data_in;
	if (addr_selector[42]&addr_selector[48])
		data_out <= r_42_48;
		if (write_en==1'b1)
			r_42_48 <= data_in;
	if (addr_selector[42]&addr_selector[49])
		data_out <= r_42_49;
		if (write_en==1'b1)
			r_42_49 <= data_in;
	if (addr_selector[42]&addr_selector[50])
		data_out <= r_42_50;
		if (write_en==1'b1)
			r_42_50 <= data_in;
	if (addr_selector[42]&addr_selector[51])
		data_out <= r_42_51;
		if (write_en==1'b1)
			r_42_51 <= data_in;
	if (addr_selector[42]&addr_selector[52])
		data_out <= r_42_52;
		if (write_en==1'b1)
			r_42_52 <= data_in;
	if (addr_selector[42]&addr_selector[53])
		data_out <= r_42_53;
		if (write_en==1'b1)
			r_42_53 <= data_in;
	if (addr_selector[42]&addr_selector[54])
		data_out <= r_42_54;
		if (write_en==1'b1)
			r_42_54 <= data_in;
	if (addr_selector[42]&addr_selector[55])
		data_out <= r_42_55;
		if (write_en==1'b1)
			r_42_55 <= data_in;
	if (addr_selector[42]&addr_selector[56])
		data_out <= r_42_56;
		if (write_en==1'b1)
			r_42_56 <= data_in;
	if (addr_selector[42]&addr_selector[57])
		data_out <= r_42_57;
		if (write_en==1'b1)
			r_42_57 <= data_in;
	if (addr_selector[42]&addr_selector[58])
		data_out <= r_42_58;
		if (write_en==1'b1)
			r_42_58 <= data_in;
	if (addr_selector[42]&addr_selector[59])
		data_out <= r_42_59;
		if (write_en==1'b1)
			r_42_59 <= data_in;
	if (addr_selector[42]&addr_selector[60])
		data_out <= r_42_60;
		if (write_en==1'b1)
			r_42_60 <= data_in;
	if (addr_selector[42]&addr_selector[61])
		data_out <= r_42_61;
		if (write_en==1'b1)
			r_42_61 <= data_in;
	if (addr_selector[42]&addr_selector[62])
		data_out <= r_42_62;
		if (write_en==1'b1)
			r_42_62 <= data_in;
	if (addr_selector[42]&addr_selector[63])
		data_out <= r_42_63;
		if (write_en==1'b1)
			r_42_63 <= data_in;
	if (addr_selector[43]&addr_selector[0])
		data_out <= r_43_0;
		if (write_en==1'b1)
			r_43_0 <= data_in;
	if (addr_selector[43]&addr_selector[1])
		data_out <= r_43_1;
		if (write_en==1'b1)
			r_43_1 <= data_in;
	if (addr_selector[43]&addr_selector[2])
		data_out <= r_43_2;
		if (write_en==1'b1)
			r_43_2 <= data_in;
	if (addr_selector[43]&addr_selector[3])
		data_out <= r_43_3;
		if (write_en==1'b1)
			r_43_3 <= data_in;
	if (addr_selector[43]&addr_selector[4])
		data_out <= r_43_4;
		if (write_en==1'b1)
			r_43_4 <= data_in;
	if (addr_selector[43]&addr_selector[5])
		data_out <= r_43_5;
		if (write_en==1'b1)
			r_43_5 <= data_in;
	if (addr_selector[43]&addr_selector[6])
		data_out <= r_43_6;
		if (write_en==1'b1)
			r_43_6 <= data_in;
	if (addr_selector[43]&addr_selector[7])
		data_out <= r_43_7;
		if (write_en==1'b1)
			r_43_7 <= data_in;
	if (addr_selector[43]&addr_selector[8])
		data_out <= r_43_8;
		if (write_en==1'b1)
			r_43_8 <= data_in;
	if (addr_selector[43]&addr_selector[9])
		data_out <= r_43_9;
		if (write_en==1'b1)
			r_43_9 <= data_in;
	if (addr_selector[43]&addr_selector[10])
		data_out <= r_43_10;
		if (write_en==1'b1)
			r_43_10 <= data_in;
	if (addr_selector[43]&addr_selector[11])
		data_out <= r_43_11;
		if (write_en==1'b1)
			r_43_11 <= data_in;
	if (addr_selector[43]&addr_selector[12])
		data_out <= r_43_12;
		if (write_en==1'b1)
			r_43_12 <= data_in;
	if (addr_selector[43]&addr_selector[13])
		data_out <= r_43_13;
		if (write_en==1'b1)
			r_43_13 <= data_in;
	if (addr_selector[43]&addr_selector[14])
		data_out <= r_43_14;
		if (write_en==1'b1)
			r_43_14 <= data_in;
	if (addr_selector[43]&addr_selector[15])
		data_out <= r_43_15;
		if (write_en==1'b1)
			r_43_15 <= data_in;
	if (addr_selector[43]&addr_selector[16])
		data_out <= r_43_16;
		if (write_en==1'b1)
			r_43_16 <= data_in;
	if (addr_selector[43]&addr_selector[17])
		data_out <= r_43_17;
		if (write_en==1'b1)
			r_43_17 <= data_in;
	if (addr_selector[43]&addr_selector[18])
		data_out <= r_43_18;
		if (write_en==1'b1)
			r_43_18 <= data_in;
	if (addr_selector[43]&addr_selector[19])
		data_out <= r_43_19;
		if (write_en==1'b1)
			r_43_19 <= data_in;
	if (addr_selector[43]&addr_selector[20])
		data_out <= r_43_20;
		if (write_en==1'b1)
			r_43_20 <= data_in;
	if (addr_selector[43]&addr_selector[21])
		data_out <= r_43_21;
		if (write_en==1'b1)
			r_43_21 <= data_in;
	if (addr_selector[43]&addr_selector[22])
		data_out <= r_43_22;
		if (write_en==1'b1)
			r_43_22 <= data_in;
	if (addr_selector[43]&addr_selector[23])
		data_out <= r_43_23;
		if (write_en==1'b1)
			r_43_23 <= data_in;
	if (addr_selector[43]&addr_selector[24])
		data_out <= r_43_24;
		if (write_en==1'b1)
			r_43_24 <= data_in;
	if (addr_selector[43]&addr_selector[25])
		data_out <= r_43_25;
		if (write_en==1'b1)
			r_43_25 <= data_in;
	if (addr_selector[43]&addr_selector[26])
		data_out <= r_43_26;
		if (write_en==1'b1)
			r_43_26 <= data_in;
	if (addr_selector[43]&addr_selector[27])
		data_out <= r_43_27;
		if (write_en==1'b1)
			r_43_27 <= data_in;
	if (addr_selector[43]&addr_selector[28])
		data_out <= r_43_28;
		if (write_en==1'b1)
			r_43_28 <= data_in;
	if (addr_selector[43]&addr_selector[29])
		data_out <= r_43_29;
		if (write_en==1'b1)
			r_43_29 <= data_in;
	if (addr_selector[43]&addr_selector[30])
		data_out <= r_43_30;
		if (write_en==1'b1)
			r_43_30 <= data_in;
	if (addr_selector[43]&addr_selector[31])
		data_out <= r_43_31;
		if (write_en==1'b1)
			r_43_31 <= data_in;
	if (addr_selector[43]&addr_selector[32])
		data_out <= r_43_32;
		if (write_en==1'b1)
			r_43_32 <= data_in;
	if (addr_selector[43]&addr_selector[33])
		data_out <= r_43_33;
		if (write_en==1'b1)
			r_43_33 <= data_in;
	if (addr_selector[43]&addr_selector[34])
		data_out <= r_43_34;
		if (write_en==1'b1)
			r_43_34 <= data_in;
	if (addr_selector[43]&addr_selector[35])
		data_out <= r_43_35;
		if (write_en==1'b1)
			r_43_35 <= data_in;
	if (addr_selector[43]&addr_selector[36])
		data_out <= r_43_36;
		if (write_en==1'b1)
			r_43_36 <= data_in;
	if (addr_selector[43]&addr_selector[37])
		data_out <= r_43_37;
		if (write_en==1'b1)
			r_43_37 <= data_in;
	if (addr_selector[43]&addr_selector[38])
		data_out <= r_43_38;
		if (write_en==1'b1)
			r_43_38 <= data_in;
	if (addr_selector[43]&addr_selector[39])
		data_out <= r_43_39;
		if (write_en==1'b1)
			r_43_39 <= data_in;
	if (addr_selector[43]&addr_selector[40])
		data_out <= r_43_40;
		if (write_en==1'b1)
			r_43_40 <= data_in;
	if (addr_selector[43]&addr_selector[41])
		data_out <= r_43_41;
		if (write_en==1'b1)
			r_43_41 <= data_in;
	if (addr_selector[43]&addr_selector[42])
		data_out <= r_43_42;
		if (write_en==1'b1)
			r_43_42 <= data_in;
	if (addr_selector[43]&addr_selector[43])
		data_out <= r_43_43;
		if (write_en==1'b1)
			r_43_43 <= data_in;
	if (addr_selector[43]&addr_selector[44])
		data_out <= r_43_44;
		if (write_en==1'b1)
			r_43_44 <= data_in;
	if (addr_selector[43]&addr_selector[45])
		data_out <= r_43_45;
		if (write_en==1'b1)
			r_43_45 <= data_in;
	if (addr_selector[43]&addr_selector[46])
		data_out <= r_43_46;
		if (write_en==1'b1)
			r_43_46 <= data_in;
	if (addr_selector[43]&addr_selector[47])
		data_out <= r_43_47;
		if (write_en==1'b1)
			r_43_47 <= data_in;
	if (addr_selector[43]&addr_selector[48])
		data_out <= r_43_48;
		if (write_en==1'b1)
			r_43_48 <= data_in;
	if (addr_selector[43]&addr_selector[49])
		data_out <= r_43_49;
		if (write_en==1'b1)
			r_43_49 <= data_in;
	if (addr_selector[43]&addr_selector[50])
		data_out <= r_43_50;
		if (write_en==1'b1)
			r_43_50 <= data_in;
	if (addr_selector[43]&addr_selector[51])
		data_out <= r_43_51;
		if (write_en==1'b1)
			r_43_51 <= data_in;
	if (addr_selector[43]&addr_selector[52])
		data_out <= r_43_52;
		if (write_en==1'b1)
			r_43_52 <= data_in;
	if (addr_selector[43]&addr_selector[53])
		data_out <= r_43_53;
		if (write_en==1'b1)
			r_43_53 <= data_in;
	if (addr_selector[43]&addr_selector[54])
		data_out <= r_43_54;
		if (write_en==1'b1)
			r_43_54 <= data_in;
	if (addr_selector[43]&addr_selector[55])
		data_out <= r_43_55;
		if (write_en==1'b1)
			r_43_55 <= data_in;
	if (addr_selector[43]&addr_selector[56])
		data_out <= r_43_56;
		if (write_en==1'b1)
			r_43_56 <= data_in;
	if (addr_selector[43]&addr_selector[57])
		data_out <= r_43_57;
		if (write_en==1'b1)
			r_43_57 <= data_in;
	if (addr_selector[43]&addr_selector[58])
		data_out <= r_43_58;
		if (write_en==1'b1)
			r_43_58 <= data_in;
	if (addr_selector[43]&addr_selector[59])
		data_out <= r_43_59;
		if (write_en==1'b1)
			r_43_59 <= data_in;
	if (addr_selector[43]&addr_selector[60])
		data_out <= r_43_60;
		if (write_en==1'b1)
			r_43_60 <= data_in;
	if (addr_selector[43]&addr_selector[61])
		data_out <= r_43_61;
		if (write_en==1'b1)
			r_43_61 <= data_in;
	if (addr_selector[43]&addr_selector[62])
		data_out <= r_43_62;
		if (write_en==1'b1)
			r_43_62 <= data_in;
	if (addr_selector[43]&addr_selector[63])
		data_out <= r_43_63;
		if (write_en==1'b1)
			r_43_63 <= data_in;
	if (addr_selector[44]&addr_selector[0])
		data_out <= r_44_0;
		if (write_en==1'b1)
			r_44_0 <= data_in;
	if (addr_selector[44]&addr_selector[1])
		data_out <= r_44_1;
		if (write_en==1'b1)
			r_44_1 <= data_in;
	if (addr_selector[44]&addr_selector[2])
		data_out <= r_44_2;
		if (write_en==1'b1)
			r_44_2 <= data_in;
	if (addr_selector[44]&addr_selector[3])
		data_out <= r_44_3;
		if (write_en==1'b1)
			r_44_3 <= data_in;
	if (addr_selector[44]&addr_selector[4])
		data_out <= r_44_4;
		if (write_en==1'b1)
			r_44_4 <= data_in;
	if (addr_selector[44]&addr_selector[5])
		data_out <= r_44_5;
		if (write_en==1'b1)
			r_44_5 <= data_in;
	if (addr_selector[44]&addr_selector[6])
		data_out <= r_44_6;
		if (write_en==1'b1)
			r_44_6 <= data_in;
	if (addr_selector[44]&addr_selector[7])
		data_out <= r_44_7;
		if (write_en==1'b1)
			r_44_7 <= data_in;
	if (addr_selector[44]&addr_selector[8])
		data_out <= r_44_8;
		if (write_en==1'b1)
			r_44_8 <= data_in;
	if (addr_selector[44]&addr_selector[9])
		data_out <= r_44_9;
		if (write_en==1'b1)
			r_44_9 <= data_in;
	if (addr_selector[44]&addr_selector[10])
		data_out <= r_44_10;
		if (write_en==1'b1)
			r_44_10 <= data_in;
	if (addr_selector[44]&addr_selector[11])
		data_out <= r_44_11;
		if (write_en==1'b1)
			r_44_11 <= data_in;
	if (addr_selector[44]&addr_selector[12])
		data_out <= r_44_12;
		if (write_en==1'b1)
			r_44_12 <= data_in;
	if (addr_selector[44]&addr_selector[13])
		data_out <= r_44_13;
		if (write_en==1'b1)
			r_44_13 <= data_in;
	if (addr_selector[44]&addr_selector[14])
		data_out <= r_44_14;
		if (write_en==1'b1)
			r_44_14 <= data_in;
	if (addr_selector[44]&addr_selector[15])
		data_out <= r_44_15;
		if (write_en==1'b1)
			r_44_15 <= data_in;
	if (addr_selector[44]&addr_selector[16])
		data_out <= r_44_16;
		if (write_en==1'b1)
			r_44_16 <= data_in;
	if (addr_selector[44]&addr_selector[17])
		data_out <= r_44_17;
		if (write_en==1'b1)
			r_44_17 <= data_in;
	if (addr_selector[44]&addr_selector[18])
		data_out <= r_44_18;
		if (write_en==1'b1)
			r_44_18 <= data_in;
	if (addr_selector[44]&addr_selector[19])
		data_out <= r_44_19;
		if (write_en==1'b1)
			r_44_19 <= data_in;
	if (addr_selector[44]&addr_selector[20])
		data_out <= r_44_20;
		if (write_en==1'b1)
			r_44_20 <= data_in;
	if (addr_selector[44]&addr_selector[21])
		data_out <= r_44_21;
		if (write_en==1'b1)
			r_44_21 <= data_in;
	if (addr_selector[44]&addr_selector[22])
		data_out <= r_44_22;
		if (write_en==1'b1)
			r_44_22 <= data_in;
	if (addr_selector[44]&addr_selector[23])
		data_out <= r_44_23;
		if (write_en==1'b1)
			r_44_23 <= data_in;
	if (addr_selector[44]&addr_selector[24])
		data_out <= r_44_24;
		if (write_en==1'b1)
			r_44_24 <= data_in;
	if (addr_selector[44]&addr_selector[25])
		data_out <= r_44_25;
		if (write_en==1'b1)
			r_44_25 <= data_in;
	if (addr_selector[44]&addr_selector[26])
		data_out <= r_44_26;
		if (write_en==1'b1)
			r_44_26 <= data_in;
	if (addr_selector[44]&addr_selector[27])
		data_out <= r_44_27;
		if (write_en==1'b1)
			r_44_27 <= data_in;
	if (addr_selector[44]&addr_selector[28])
		data_out <= r_44_28;
		if (write_en==1'b1)
			r_44_28 <= data_in;
	if (addr_selector[44]&addr_selector[29])
		data_out <= r_44_29;
		if (write_en==1'b1)
			r_44_29 <= data_in;
	if (addr_selector[44]&addr_selector[30])
		data_out <= r_44_30;
		if (write_en==1'b1)
			r_44_30 <= data_in;
	if (addr_selector[44]&addr_selector[31])
		data_out <= r_44_31;
		if (write_en==1'b1)
			r_44_31 <= data_in;
	if (addr_selector[44]&addr_selector[32])
		data_out <= r_44_32;
		if (write_en==1'b1)
			r_44_32 <= data_in;
	if (addr_selector[44]&addr_selector[33])
		data_out <= r_44_33;
		if (write_en==1'b1)
			r_44_33 <= data_in;
	if (addr_selector[44]&addr_selector[34])
		data_out <= r_44_34;
		if (write_en==1'b1)
			r_44_34 <= data_in;
	if (addr_selector[44]&addr_selector[35])
		data_out <= r_44_35;
		if (write_en==1'b1)
			r_44_35 <= data_in;
	if (addr_selector[44]&addr_selector[36])
		data_out <= r_44_36;
		if (write_en==1'b1)
			r_44_36 <= data_in;
	if (addr_selector[44]&addr_selector[37])
		data_out <= r_44_37;
		if (write_en==1'b1)
			r_44_37 <= data_in;
	if (addr_selector[44]&addr_selector[38])
		data_out <= r_44_38;
		if (write_en==1'b1)
			r_44_38 <= data_in;
	if (addr_selector[44]&addr_selector[39])
		data_out <= r_44_39;
		if (write_en==1'b1)
			r_44_39 <= data_in;
	if (addr_selector[44]&addr_selector[40])
		data_out <= r_44_40;
		if (write_en==1'b1)
			r_44_40 <= data_in;
	if (addr_selector[44]&addr_selector[41])
		data_out <= r_44_41;
		if (write_en==1'b1)
			r_44_41 <= data_in;
	if (addr_selector[44]&addr_selector[42])
		data_out <= r_44_42;
		if (write_en==1'b1)
			r_44_42 <= data_in;
	if (addr_selector[44]&addr_selector[43])
		data_out <= r_44_43;
		if (write_en==1'b1)
			r_44_43 <= data_in;
	if (addr_selector[44]&addr_selector[44])
		data_out <= r_44_44;
		if (write_en==1'b1)
			r_44_44 <= data_in;
	if (addr_selector[44]&addr_selector[45])
		data_out <= r_44_45;
		if (write_en==1'b1)
			r_44_45 <= data_in;
	if (addr_selector[44]&addr_selector[46])
		data_out <= r_44_46;
		if (write_en==1'b1)
			r_44_46 <= data_in;
	if (addr_selector[44]&addr_selector[47])
		data_out <= r_44_47;
		if (write_en==1'b1)
			r_44_47 <= data_in;
	if (addr_selector[44]&addr_selector[48])
		data_out <= r_44_48;
		if (write_en==1'b1)
			r_44_48 <= data_in;
	if (addr_selector[44]&addr_selector[49])
		data_out <= r_44_49;
		if (write_en==1'b1)
			r_44_49 <= data_in;
	if (addr_selector[44]&addr_selector[50])
		data_out <= r_44_50;
		if (write_en==1'b1)
			r_44_50 <= data_in;
	if (addr_selector[44]&addr_selector[51])
		data_out <= r_44_51;
		if (write_en==1'b1)
			r_44_51 <= data_in;
	if (addr_selector[44]&addr_selector[52])
		data_out <= r_44_52;
		if (write_en==1'b1)
			r_44_52 <= data_in;
	if (addr_selector[44]&addr_selector[53])
		data_out <= r_44_53;
		if (write_en==1'b1)
			r_44_53 <= data_in;
	if (addr_selector[44]&addr_selector[54])
		data_out <= r_44_54;
		if (write_en==1'b1)
			r_44_54 <= data_in;
	if (addr_selector[44]&addr_selector[55])
		data_out <= r_44_55;
		if (write_en==1'b1)
			r_44_55 <= data_in;
	if (addr_selector[44]&addr_selector[56])
		data_out <= r_44_56;
		if (write_en==1'b1)
			r_44_56 <= data_in;
	if (addr_selector[44]&addr_selector[57])
		data_out <= r_44_57;
		if (write_en==1'b1)
			r_44_57 <= data_in;
	if (addr_selector[44]&addr_selector[58])
		data_out <= r_44_58;
		if (write_en==1'b1)
			r_44_58 <= data_in;
	if (addr_selector[44]&addr_selector[59])
		data_out <= r_44_59;
		if (write_en==1'b1)
			r_44_59 <= data_in;
	if (addr_selector[44]&addr_selector[60])
		data_out <= r_44_60;
		if (write_en==1'b1)
			r_44_60 <= data_in;
	if (addr_selector[44]&addr_selector[61])
		data_out <= r_44_61;
		if (write_en==1'b1)
			r_44_61 <= data_in;
	if (addr_selector[44]&addr_selector[62])
		data_out <= r_44_62;
		if (write_en==1'b1)
			r_44_62 <= data_in;
	if (addr_selector[44]&addr_selector[63])
		data_out <= r_44_63;
		if (write_en==1'b1)
			r_44_63 <= data_in;
	if (addr_selector[45]&addr_selector[0])
		data_out <= r_45_0;
		if (write_en==1'b1)
			r_45_0 <= data_in;
	if (addr_selector[45]&addr_selector[1])
		data_out <= r_45_1;
		if (write_en==1'b1)
			r_45_1 <= data_in;
	if (addr_selector[45]&addr_selector[2])
		data_out <= r_45_2;
		if (write_en==1'b1)
			r_45_2 <= data_in;
	if (addr_selector[45]&addr_selector[3])
		data_out <= r_45_3;
		if (write_en==1'b1)
			r_45_3 <= data_in;
	if (addr_selector[45]&addr_selector[4])
		data_out <= r_45_4;
		if (write_en==1'b1)
			r_45_4 <= data_in;
	if (addr_selector[45]&addr_selector[5])
		data_out <= r_45_5;
		if (write_en==1'b1)
			r_45_5 <= data_in;
	if (addr_selector[45]&addr_selector[6])
		data_out <= r_45_6;
		if (write_en==1'b1)
			r_45_6 <= data_in;
	if (addr_selector[45]&addr_selector[7])
		data_out <= r_45_7;
		if (write_en==1'b1)
			r_45_7 <= data_in;
	if (addr_selector[45]&addr_selector[8])
		data_out <= r_45_8;
		if (write_en==1'b1)
			r_45_8 <= data_in;
	if (addr_selector[45]&addr_selector[9])
		data_out <= r_45_9;
		if (write_en==1'b1)
			r_45_9 <= data_in;
	if (addr_selector[45]&addr_selector[10])
		data_out <= r_45_10;
		if (write_en==1'b1)
			r_45_10 <= data_in;
	if (addr_selector[45]&addr_selector[11])
		data_out <= r_45_11;
		if (write_en==1'b1)
			r_45_11 <= data_in;
	if (addr_selector[45]&addr_selector[12])
		data_out <= r_45_12;
		if (write_en==1'b1)
			r_45_12 <= data_in;
	if (addr_selector[45]&addr_selector[13])
		data_out <= r_45_13;
		if (write_en==1'b1)
			r_45_13 <= data_in;
	if (addr_selector[45]&addr_selector[14])
		data_out <= r_45_14;
		if (write_en==1'b1)
			r_45_14 <= data_in;
	if (addr_selector[45]&addr_selector[15])
		data_out <= r_45_15;
		if (write_en==1'b1)
			r_45_15 <= data_in;
	if (addr_selector[45]&addr_selector[16])
		data_out <= r_45_16;
		if (write_en==1'b1)
			r_45_16 <= data_in;
	if (addr_selector[45]&addr_selector[17])
		data_out <= r_45_17;
		if (write_en==1'b1)
			r_45_17 <= data_in;
	if (addr_selector[45]&addr_selector[18])
		data_out <= r_45_18;
		if (write_en==1'b1)
			r_45_18 <= data_in;
	if (addr_selector[45]&addr_selector[19])
		data_out <= r_45_19;
		if (write_en==1'b1)
			r_45_19 <= data_in;
	if (addr_selector[45]&addr_selector[20])
		data_out <= r_45_20;
		if (write_en==1'b1)
			r_45_20 <= data_in;
	if (addr_selector[45]&addr_selector[21])
		data_out <= r_45_21;
		if (write_en==1'b1)
			r_45_21 <= data_in;
	if (addr_selector[45]&addr_selector[22])
		data_out <= r_45_22;
		if (write_en==1'b1)
			r_45_22 <= data_in;
	if (addr_selector[45]&addr_selector[23])
		data_out <= r_45_23;
		if (write_en==1'b1)
			r_45_23 <= data_in;
	if (addr_selector[45]&addr_selector[24])
		data_out <= r_45_24;
		if (write_en==1'b1)
			r_45_24 <= data_in;
	if (addr_selector[45]&addr_selector[25])
		data_out <= r_45_25;
		if (write_en==1'b1)
			r_45_25 <= data_in;
	if (addr_selector[45]&addr_selector[26])
		data_out <= r_45_26;
		if (write_en==1'b1)
			r_45_26 <= data_in;
	if (addr_selector[45]&addr_selector[27])
		data_out <= r_45_27;
		if (write_en==1'b1)
			r_45_27 <= data_in;
	if (addr_selector[45]&addr_selector[28])
		data_out <= r_45_28;
		if (write_en==1'b1)
			r_45_28 <= data_in;
	if (addr_selector[45]&addr_selector[29])
		data_out <= r_45_29;
		if (write_en==1'b1)
			r_45_29 <= data_in;
	if (addr_selector[45]&addr_selector[30])
		data_out <= r_45_30;
		if (write_en==1'b1)
			r_45_30 <= data_in;
	if (addr_selector[45]&addr_selector[31])
		data_out <= r_45_31;
		if (write_en==1'b1)
			r_45_31 <= data_in;
	if (addr_selector[45]&addr_selector[32])
		data_out <= r_45_32;
		if (write_en==1'b1)
			r_45_32 <= data_in;
	if (addr_selector[45]&addr_selector[33])
		data_out <= r_45_33;
		if (write_en==1'b1)
			r_45_33 <= data_in;
	if (addr_selector[45]&addr_selector[34])
		data_out <= r_45_34;
		if (write_en==1'b1)
			r_45_34 <= data_in;
	if (addr_selector[45]&addr_selector[35])
		data_out <= r_45_35;
		if (write_en==1'b1)
			r_45_35 <= data_in;
	if (addr_selector[45]&addr_selector[36])
		data_out <= r_45_36;
		if (write_en==1'b1)
			r_45_36 <= data_in;
	if (addr_selector[45]&addr_selector[37])
		data_out <= r_45_37;
		if (write_en==1'b1)
			r_45_37 <= data_in;
	if (addr_selector[45]&addr_selector[38])
		data_out <= r_45_38;
		if (write_en==1'b1)
			r_45_38 <= data_in;
	if (addr_selector[45]&addr_selector[39])
		data_out <= r_45_39;
		if (write_en==1'b1)
			r_45_39 <= data_in;
	if (addr_selector[45]&addr_selector[40])
		data_out <= r_45_40;
		if (write_en==1'b1)
			r_45_40 <= data_in;
	if (addr_selector[45]&addr_selector[41])
		data_out <= r_45_41;
		if (write_en==1'b1)
			r_45_41 <= data_in;
	if (addr_selector[45]&addr_selector[42])
		data_out <= r_45_42;
		if (write_en==1'b1)
			r_45_42 <= data_in;
	if (addr_selector[45]&addr_selector[43])
		data_out <= r_45_43;
		if (write_en==1'b1)
			r_45_43 <= data_in;
	if (addr_selector[45]&addr_selector[44])
		data_out <= r_45_44;
		if (write_en==1'b1)
			r_45_44 <= data_in;
	if (addr_selector[45]&addr_selector[45])
		data_out <= r_45_45;
		if (write_en==1'b1)
			r_45_45 <= data_in;
	if (addr_selector[45]&addr_selector[46])
		data_out <= r_45_46;
		if (write_en==1'b1)
			r_45_46 <= data_in;
	if (addr_selector[45]&addr_selector[47])
		data_out <= r_45_47;
		if (write_en==1'b1)
			r_45_47 <= data_in;
	if (addr_selector[45]&addr_selector[48])
		data_out <= r_45_48;
		if (write_en==1'b1)
			r_45_48 <= data_in;
	if (addr_selector[45]&addr_selector[49])
		data_out <= r_45_49;
		if (write_en==1'b1)
			r_45_49 <= data_in;
	if (addr_selector[45]&addr_selector[50])
		data_out <= r_45_50;
		if (write_en==1'b1)
			r_45_50 <= data_in;
	if (addr_selector[45]&addr_selector[51])
		data_out <= r_45_51;
		if (write_en==1'b1)
			r_45_51 <= data_in;
	if (addr_selector[45]&addr_selector[52])
		data_out <= r_45_52;
		if (write_en==1'b1)
			r_45_52 <= data_in;
	if (addr_selector[45]&addr_selector[53])
		data_out <= r_45_53;
		if (write_en==1'b1)
			r_45_53 <= data_in;
	if (addr_selector[45]&addr_selector[54])
		data_out <= r_45_54;
		if (write_en==1'b1)
			r_45_54 <= data_in;
	if (addr_selector[45]&addr_selector[55])
		data_out <= r_45_55;
		if (write_en==1'b1)
			r_45_55 <= data_in;
	if (addr_selector[45]&addr_selector[56])
		data_out <= r_45_56;
		if (write_en==1'b1)
			r_45_56 <= data_in;
	if (addr_selector[45]&addr_selector[57])
		data_out <= r_45_57;
		if (write_en==1'b1)
			r_45_57 <= data_in;
	if (addr_selector[45]&addr_selector[58])
		data_out <= r_45_58;
		if (write_en==1'b1)
			r_45_58 <= data_in;
	if (addr_selector[45]&addr_selector[59])
		data_out <= r_45_59;
		if (write_en==1'b1)
			r_45_59 <= data_in;
	if (addr_selector[45]&addr_selector[60])
		data_out <= r_45_60;
		if (write_en==1'b1)
			r_45_60 <= data_in;
	if (addr_selector[45]&addr_selector[61])
		data_out <= r_45_61;
		if (write_en==1'b1)
			r_45_61 <= data_in;
	if (addr_selector[45]&addr_selector[62])
		data_out <= r_45_62;
		if (write_en==1'b1)
			r_45_62 <= data_in;
	if (addr_selector[45]&addr_selector[63])
		data_out <= r_45_63;
		if (write_en==1'b1)
			r_45_63 <= data_in;
	if (addr_selector[46]&addr_selector[0])
		data_out <= r_46_0;
		if (write_en==1'b1)
			r_46_0 <= data_in;
	if (addr_selector[46]&addr_selector[1])
		data_out <= r_46_1;
		if (write_en==1'b1)
			r_46_1 <= data_in;
	if (addr_selector[46]&addr_selector[2])
		data_out <= r_46_2;
		if (write_en==1'b1)
			r_46_2 <= data_in;
	if (addr_selector[46]&addr_selector[3])
		data_out <= r_46_3;
		if (write_en==1'b1)
			r_46_3 <= data_in;
	if (addr_selector[46]&addr_selector[4])
		data_out <= r_46_4;
		if (write_en==1'b1)
			r_46_4 <= data_in;
	if (addr_selector[46]&addr_selector[5])
		data_out <= r_46_5;
		if (write_en==1'b1)
			r_46_5 <= data_in;
	if (addr_selector[46]&addr_selector[6])
		data_out <= r_46_6;
		if (write_en==1'b1)
			r_46_6 <= data_in;
	if (addr_selector[46]&addr_selector[7])
		data_out <= r_46_7;
		if (write_en==1'b1)
			r_46_7 <= data_in;
	if (addr_selector[46]&addr_selector[8])
		data_out <= r_46_8;
		if (write_en==1'b1)
			r_46_8 <= data_in;
	if (addr_selector[46]&addr_selector[9])
		data_out <= r_46_9;
		if (write_en==1'b1)
			r_46_9 <= data_in;
	if (addr_selector[46]&addr_selector[10])
		data_out <= r_46_10;
		if (write_en==1'b1)
			r_46_10 <= data_in;
	if (addr_selector[46]&addr_selector[11])
		data_out <= r_46_11;
		if (write_en==1'b1)
			r_46_11 <= data_in;
	if (addr_selector[46]&addr_selector[12])
		data_out <= r_46_12;
		if (write_en==1'b1)
			r_46_12 <= data_in;
	if (addr_selector[46]&addr_selector[13])
		data_out <= r_46_13;
		if (write_en==1'b1)
			r_46_13 <= data_in;
	if (addr_selector[46]&addr_selector[14])
		data_out <= r_46_14;
		if (write_en==1'b1)
			r_46_14 <= data_in;
	if (addr_selector[46]&addr_selector[15])
		data_out <= r_46_15;
		if (write_en==1'b1)
			r_46_15 <= data_in;
	if (addr_selector[46]&addr_selector[16])
		data_out <= r_46_16;
		if (write_en==1'b1)
			r_46_16 <= data_in;
	if (addr_selector[46]&addr_selector[17])
		data_out <= r_46_17;
		if (write_en==1'b1)
			r_46_17 <= data_in;
	if (addr_selector[46]&addr_selector[18])
		data_out <= r_46_18;
		if (write_en==1'b1)
			r_46_18 <= data_in;
	if (addr_selector[46]&addr_selector[19])
		data_out <= r_46_19;
		if (write_en==1'b1)
			r_46_19 <= data_in;
	if (addr_selector[46]&addr_selector[20])
		data_out <= r_46_20;
		if (write_en==1'b1)
			r_46_20 <= data_in;
	if (addr_selector[46]&addr_selector[21])
		data_out <= r_46_21;
		if (write_en==1'b1)
			r_46_21 <= data_in;
	if (addr_selector[46]&addr_selector[22])
		data_out <= r_46_22;
		if (write_en==1'b1)
			r_46_22 <= data_in;
	if (addr_selector[46]&addr_selector[23])
		data_out <= r_46_23;
		if (write_en==1'b1)
			r_46_23 <= data_in;
	if (addr_selector[46]&addr_selector[24])
		data_out <= r_46_24;
		if (write_en==1'b1)
			r_46_24 <= data_in;
	if (addr_selector[46]&addr_selector[25])
		data_out <= r_46_25;
		if (write_en==1'b1)
			r_46_25 <= data_in;
	if (addr_selector[46]&addr_selector[26])
		data_out <= r_46_26;
		if (write_en==1'b1)
			r_46_26 <= data_in;
	if (addr_selector[46]&addr_selector[27])
		data_out <= r_46_27;
		if (write_en==1'b1)
			r_46_27 <= data_in;
	if (addr_selector[46]&addr_selector[28])
		data_out <= r_46_28;
		if (write_en==1'b1)
			r_46_28 <= data_in;
	if (addr_selector[46]&addr_selector[29])
		data_out <= r_46_29;
		if (write_en==1'b1)
			r_46_29 <= data_in;
	if (addr_selector[46]&addr_selector[30])
		data_out <= r_46_30;
		if (write_en==1'b1)
			r_46_30 <= data_in;
	if (addr_selector[46]&addr_selector[31])
		data_out <= r_46_31;
		if (write_en==1'b1)
			r_46_31 <= data_in;
	if (addr_selector[46]&addr_selector[32])
		data_out <= r_46_32;
		if (write_en==1'b1)
			r_46_32 <= data_in;
	if (addr_selector[46]&addr_selector[33])
		data_out <= r_46_33;
		if (write_en==1'b1)
			r_46_33 <= data_in;
	if (addr_selector[46]&addr_selector[34])
		data_out <= r_46_34;
		if (write_en==1'b1)
			r_46_34 <= data_in;
	if (addr_selector[46]&addr_selector[35])
		data_out <= r_46_35;
		if (write_en==1'b1)
			r_46_35 <= data_in;
	if (addr_selector[46]&addr_selector[36])
		data_out <= r_46_36;
		if (write_en==1'b1)
			r_46_36 <= data_in;
	if (addr_selector[46]&addr_selector[37])
		data_out <= r_46_37;
		if (write_en==1'b1)
			r_46_37 <= data_in;
	if (addr_selector[46]&addr_selector[38])
		data_out <= r_46_38;
		if (write_en==1'b1)
			r_46_38 <= data_in;
	if (addr_selector[46]&addr_selector[39])
		data_out <= r_46_39;
		if (write_en==1'b1)
			r_46_39 <= data_in;
	if (addr_selector[46]&addr_selector[40])
		data_out <= r_46_40;
		if (write_en==1'b1)
			r_46_40 <= data_in;
	if (addr_selector[46]&addr_selector[41])
		data_out <= r_46_41;
		if (write_en==1'b1)
			r_46_41 <= data_in;
	if (addr_selector[46]&addr_selector[42])
		data_out <= r_46_42;
		if (write_en==1'b1)
			r_46_42 <= data_in;
	if (addr_selector[46]&addr_selector[43])
		data_out <= r_46_43;
		if (write_en==1'b1)
			r_46_43 <= data_in;
	if (addr_selector[46]&addr_selector[44])
		data_out <= r_46_44;
		if (write_en==1'b1)
			r_46_44 <= data_in;
	if (addr_selector[46]&addr_selector[45])
		data_out <= r_46_45;
		if (write_en==1'b1)
			r_46_45 <= data_in;
	if (addr_selector[46]&addr_selector[46])
		data_out <= r_46_46;
		if (write_en==1'b1)
			r_46_46 <= data_in;
	if (addr_selector[46]&addr_selector[47])
		data_out <= r_46_47;
		if (write_en==1'b1)
			r_46_47 <= data_in;
	if (addr_selector[46]&addr_selector[48])
		data_out <= r_46_48;
		if (write_en==1'b1)
			r_46_48 <= data_in;
	if (addr_selector[46]&addr_selector[49])
		data_out <= r_46_49;
		if (write_en==1'b1)
			r_46_49 <= data_in;
	if (addr_selector[46]&addr_selector[50])
		data_out <= r_46_50;
		if (write_en==1'b1)
			r_46_50 <= data_in;
	if (addr_selector[46]&addr_selector[51])
		data_out <= r_46_51;
		if (write_en==1'b1)
			r_46_51 <= data_in;
	if (addr_selector[46]&addr_selector[52])
		data_out <= r_46_52;
		if (write_en==1'b1)
			r_46_52 <= data_in;
	if (addr_selector[46]&addr_selector[53])
		data_out <= r_46_53;
		if (write_en==1'b1)
			r_46_53 <= data_in;
	if (addr_selector[46]&addr_selector[54])
		data_out <= r_46_54;
		if (write_en==1'b1)
			r_46_54 <= data_in;
	if (addr_selector[46]&addr_selector[55])
		data_out <= r_46_55;
		if (write_en==1'b1)
			r_46_55 <= data_in;
	if (addr_selector[46]&addr_selector[56])
		data_out <= r_46_56;
		if (write_en==1'b1)
			r_46_56 <= data_in;
	if (addr_selector[46]&addr_selector[57])
		data_out <= r_46_57;
		if (write_en==1'b1)
			r_46_57 <= data_in;
	if (addr_selector[46]&addr_selector[58])
		data_out <= r_46_58;
		if (write_en==1'b1)
			r_46_58 <= data_in;
	if (addr_selector[46]&addr_selector[59])
		data_out <= r_46_59;
		if (write_en==1'b1)
			r_46_59 <= data_in;
	if (addr_selector[46]&addr_selector[60])
		data_out <= r_46_60;
		if (write_en==1'b1)
			r_46_60 <= data_in;
	if (addr_selector[46]&addr_selector[61])
		data_out <= r_46_61;
		if (write_en==1'b1)
			r_46_61 <= data_in;
	if (addr_selector[46]&addr_selector[62])
		data_out <= r_46_62;
		if (write_en==1'b1)
			r_46_62 <= data_in;
	if (addr_selector[46]&addr_selector[63])
		data_out <= r_46_63;
		if (write_en==1'b1)
			r_46_63 <= data_in;
	if (addr_selector[47]&addr_selector[0])
		data_out <= r_47_0;
		if (write_en==1'b1)
			r_47_0 <= data_in;
	if (addr_selector[47]&addr_selector[1])
		data_out <= r_47_1;
		if (write_en==1'b1)
			r_47_1 <= data_in;
	if (addr_selector[47]&addr_selector[2])
		data_out <= r_47_2;
		if (write_en==1'b1)
			r_47_2 <= data_in;
	if (addr_selector[47]&addr_selector[3])
		data_out <= r_47_3;
		if (write_en==1'b1)
			r_47_3 <= data_in;
	if (addr_selector[47]&addr_selector[4])
		data_out <= r_47_4;
		if (write_en==1'b1)
			r_47_4 <= data_in;
	if (addr_selector[47]&addr_selector[5])
		data_out <= r_47_5;
		if (write_en==1'b1)
			r_47_5 <= data_in;
	if (addr_selector[47]&addr_selector[6])
		data_out <= r_47_6;
		if (write_en==1'b1)
			r_47_6 <= data_in;
	if (addr_selector[47]&addr_selector[7])
		data_out <= r_47_7;
		if (write_en==1'b1)
			r_47_7 <= data_in;
	if (addr_selector[47]&addr_selector[8])
		data_out <= r_47_8;
		if (write_en==1'b1)
			r_47_8 <= data_in;
	if (addr_selector[47]&addr_selector[9])
		data_out <= r_47_9;
		if (write_en==1'b1)
			r_47_9 <= data_in;
	if (addr_selector[47]&addr_selector[10])
		data_out <= r_47_10;
		if (write_en==1'b1)
			r_47_10 <= data_in;
	if (addr_selector[47]&addr_selector[11])
		data_out <= r_47_11;
		if (write_en==1'b1)
			r_47_11 <= data_in;
	if (addr_selector[47]&addr_selector[12])
		data_out <= r_47_12;
		if (write_en==1'b1)
			r_47_12 <= data_in;
	if (addr_selector[47]&addr_selector[13])
		data_out <= r_47_13;
		if (write_en==1'b1)
			r_47_13 <= data_in;
	if (addr_selector[47]&addr_selector[14])
		data_out <= r_47_14;
		if (write_en==1'b1)
			r_47_14 <= data_in;
	if (addr_selector[47]&addr_selector[15])
		data_out <= r_47_15;
		if (write_en==1'b1)
			r_47_15 <= data_in;
	if (addr_selector[47]&addr_selector[16])
		data_out <= r_47_16;
		if (write_en==1'b1)
			r_47_16 <= data_in;
	if (addr_selector[47]&addr_selector[17])
		data_out <= r_47_17;
		if (write_en==1'b1)
			r_47_17 <= data_in;
	if (addr_selector[47]&addr_selector[18])
		data_out <= r_47_18;
		if (write_en==1'b1)
			r_47_18 <= data_in;
	if (addr_selector[47]&addr_selector[19])
		data_out <= r_47_19;
		if (write_en==1'b1)
			r_47_19 <= data_in;
	if (addr_selector[47]&addr_selector[20])
		data_out <= r_47_20;
		if (write_en==1'b1)
			r_47_20 <= data_in;
	if (addr_selector[47]&addr_selector[21])
		data_out <= r_47_21;
		if (write_en==1'b1)
			r_47_21 <= data_in;
	if (addr_selector[47]&addr_selector[22])
		data_out <= r_47_22;
		if (write_en==1'b1)
			r_47_22 <= data_in;
	if (addr_selector[47]&addr_selector[23])
		data_out <= r_47_23;
		if (write_en==1'b1)
			r_47_23 <= data_in;
	if (addr_selector[47]&addr_selector[24])
		data_out <= r_47_24;
		if (write_en==1'b1)
			r_47_24 <= data_in;
	if (addr_selector[47]&addr_selector[25])
		data_out <= r_47_25;
		if (write_en==1'b1)
			r_47_25 <= data_in;
	if (addr_selector[47]&addr_selector[26])
		data_out <= r_47_26;
		if (write_en==1'b1)
			r_47_26 <= data_in;
	if (addr_selector[47]&addr_selector[27])
		data_out <= r_47_27;
		if (write_en==1'b1)
			r_47_27 <= data_in;
	if (addr_selector[47]&addr_selector[28])
		data_out <= r_47_28;
		if (write_en==1'b1)
			r_47_28 <= data_in;
	if (addr_selector[47]&addr_selector[29])
		data_out <= r_47_29;
		if (write_en==1'b1)
			r_47_29 <= data_in;
	if (addr_selector[47]&addr_selector[30])
		data_out <= r_47_30;
		if (write_en==1'b1)
			r_47_30 <= data_in;
	if (addr_selector[47]&addr_selector[31])
		data_out <= r_47_31;
		if (write_en==1'b1)
			r_47_31 <= data_in;
	if (addr_selector[47]&addr_selector[32])
		data_out <= r_47_32;
		if (write_en==1'b1)
			r_47_32 <= data_in;
	if (addr_selector[47]&addr_selector[33])
		data_out <= r_47_33;
		if (write_en==1'b1)
			r_47_33 <= data_in;
	if (addr_selector[47]&addr_selector[34])
		data_out <= r_47_34;
		if (write_en==1'b1)
			r_47_34 <= data_in;
	if (addr_selector[47]&addr_selector[35])
		data_out <= r_47_35;
		if (write_en==1'b1)
			r_47_35 <= data_in;
	if (addr_selector[47]&addr_selector[36])
		data_out <= r_47_36;
		if (write_en==1'b1)
			r_47_36 <= data_in;
	if (addr_selector[47]&addr_selector[37])
		data_out <= r_47_37;
		if (write_en==1'b1)
			r_47_37 <= data_in;
	if (addr_selector[47]&addr_selector[38])
		data_out <= r_47_38;
		if (write_en==1'b1)
			r_47_38 <= data_in;
	if (addr_selector[47]&addr_selector[39])
		data_out <= r_47_39;
		if (write_en==1'b1)
			r_47_39 <= data_in;
	if (addr_selector[47]&addr_selector[40])
		data_out <= r_47_40;
		if (write_en==1'b1)
			r_47_40 <= data_in;
	if (addr_selector[47]&addr_selector[41])
		data_out <= r_47_41;
		if (write_en==1'b1)
			r_47_41 <= data_in;
	if (addr_selector[47]&addr_selector[42])
		data_out <= r_47_42;
		if (write_en==1'b1)
			r_47_42 <= data_in;
	if (addr_selector[47]&addr_selector[43])
		data_out <= r_47_43;
		if (write_en==1'b1)
			r_47_43 <= data_in;
	if (addr_selector[47]&addr_selector[44])
		data_out <= r_47_44;
		if (write_en==1'b1)
			r_47_44 <= data_in;
	if (addr_selector[47]&addr_selector[45])
		data_out <= r_47_45;
		if (write_en==1'b1)
			r_47_45 <= data_in;
	if (addr_selector[47]&addr_selector[46])
		data_out <= r_47_46;
		if (write_en==1'b1)
			r_47_46 <= data_in;
	if (addr_selector[47]&addr_selector[47])
		data_out <= r_47_47;
		if (write_en==1'b1)
			r_47_47 <= data_in;
	if (addr_selector[47]&addr_selector[48])
		data_out <= r_47_48;
		if (write_en==1'b1)
			r_47_48 <= data_in;
	if (addr_selector[47]&addr_selector[49])
		data_out <= r_47_49;
		if (write_en==1'b1)
			r_47_49 <= data_in;
	if (addr_selector[47]&addr_selector[50])
		data_out <= r_47_50;
		if (write_en==1'b1)
			r_47_50 <= data_in;
	if (addr_selector[47]&addr_selector[51])
		data_out <= r_47_51;
		if (write_en==1'b1)
			r_47_51 <= data_in;
	if (addr_selector[47]&addr_selector[52])
		data_out <= r_47_52;
		if (write_en==1'b1)
			r_47_52 <= data_in;
	if (addr_selector[47]&addr_selector[53])
		data_out <= r_47_53;
		if (write_en==1'b1)
			r_47_53 <= data_in;
	if (addr_selector[47]&addr_selector[54])
		data_out <= r_47_54;
		if (write_en==1'b1)
			r_47_54 <= data_in;
	if (addr_selector[47]&addr_selector[55])
		data_out <= r_47_55;
		if (write_en==1'b1)
			r_47_55 <= data_in;
	if (addr_selector[47]&addr_selector[56])
		data_out <= r_47_56;
		if (write_en==1'b1)
			r_47_56 <= data_in;
	if (addr_selector[47]&addr_selector[57])
		data_out <= r_47_57;
		if (write_en==1'b1)
			r_47_57 <= data_in;
	if (addr_selector[47]&addr_selector[58])
		data_out <= r_47_58;
		if (write_en==1'b1)
			r_47_58 <= data_in;
	if (addr_selector[47]&addr_selector[59])
		data_out <= r_47_59;
		if (write_en==1'b1)
			r_47_59 <= data_in;
	if (addr_selector[47]&addr_selector[60])
		data_out <= r_47_60;
		if (write_en==1'b1)
			r_47_60 <= data_in;
	if (addr_selector[47]&addr_selector[61])
		data_out <= r_47_61;
		if (write_en==1'b1)
			r_47_61 <= data_in;
	if (addr_selector[47]&addr_selector[62])
		data_out <= r_47_62;
		if (write_en==1'b1)
			r_47_62 <= data_in;
	if (addr_selector[47]&addr_selector[63])
		data_out <= r_47_63;
		if (write_en==1'b1)
			r_47_63 <= data_in;
	if (addr_selector[48]&addr_selector[0])
		data_out <= r_48_0;
		if (write_en==1'b1)
			r_48_0 <= data_in;
	if (addr_selector[48]&addr_selector[1])
		data_out <= r_48_1;
		if (write_en==1'b1)
			r_48_1 <= data_in;
	if (addr_selector[48]&addr_selector[2])
		data_out <= r_48_2;
		if (write_en==1'b1)
			r_48_2 <= data_in;
	if (addr_selector[48]&addr_selector[3])
		data_out <= r_48_3;
		if (write_en==1'b1)
			r_48_3 <= data_in;
	if (addr_selector[48]&addr_selector[4])
		data_out <= r_48_4;
		if (write_en==1'b1)
			r_48_4 <= data_in;
	if (addr_selector[48]&addr_selector[5])
		data_out <= r_48_5;
		if (write_en==1'b1)
			r_48_5 <= data_in;
	if (addr_selector[48]&addr_selector[6])
		data_out <= r_48_6;
		if (write_en==1'b1)
			r_48_6 <= data_in;
	if (addr_selector[48]&addr_selector[7])
		data_out <= r_48_7;
		if (write_en==1'b1)
			r_48_7 <= data_in;
	if (addr_selector[48]&addr_selector[8])
		data_out <= r_48_8;
		if (write_en==1'b1)
			r_48_8 <= data_in;
	if (addr_selector[48]&addr_selector[9])
		data_out <= r_48_9;
		if (write_en==1'b1)
			r_48_9 <= data_in;
	if (addr_selector[48]&addr_selector[10])
		data_out <= r_48_10;
		if (write_en==1'b1)
			r_48_10 <= data_in;
	if (addr_selector[48]&addr_selector[11])
		data_out <= r_48_11;
		if (write_en==1'b1)
			r_48_11 <= data_in;
	if (addr_selector[48]&addr_selector[12])
		data_out <= r_48_12;
		if (write_en==1'b1)
			r_48_12 <= data_in;
	if (addr_selector[48]&addr_selector[13])
		data_out <= r_48_13;
		if (write_en==1'b1)
			r_48_13 <= data_in;
	if (addr_selector[48]&addr_selector[14])
		data_out <= r_48_14;
		if (write_en==1'b1)
			r_48_14 <= data_in;
	if (addr_selector[48]&addr_selector[15])
		data_out <= r_48_15;
		if (write_en==1'b1)
			r_48_15 <= data_in;
	if (addr_selector[48]&addr_selector[16])
		data_out <= r_48_16;
		if (write_en==1'b1)
			r_48_16 <= data_in;
	if (addr_selector[48]&addr_selector[17])
		data_out <= r_48_17;
		if (write_en==1'b1)
			r_48_17 <= data_in;
	if (addr_selector[48]&addr_selector[18])
		data_out <= r_48_18;
		if (write_en==1'b1)
			r_48_18 <= data_in;
	if (addr_selector[48]&addr_selector[19])
		data_out <= r_48_19;
		if (write_en==1'b1)
			r_48_19 <= data_in;
	if (addr_selector[48]&addr_selector[20])
		data_out <= r_48_20;
		if (write_en==1'b1)
			r_48_20 <= data_in;
	if (addr_selector[48]&addr_selector[21])
		data_out <= r_48_21;
		if (write_en==1'b1)
			r_48_21 <= data_in;
	if (addr_selector[48]&addr_selector[22])
		data_out <= r_48_22;
		if (write_en==1'b1)
			r_48_22 <= data_in;
	if (addr_selector[48]&addr_selector[23])
		data_out <= r_48_23;
		if (write_en==1'b1)
			r_48_23 <= data_in;
	if (addr_selector[48]&addr_selector[24])
		data_out <= r_48_24;
		if (write_en==1'b1)
			r_48_24 <= data_in;
	if (addr_selector[48]&addr_selector[25])
		data_out <= r_48_25;
		if (write_en==1'b1)
			r_48_25 <= data_in;
	if (addr_selector[48]&addr_selector[26])
		data_out <= r_48_26;
		if (write_en==1'b1)
			r_48_26 <= data_in;
	if (addr_selector[48]&addr_selector[27])
		data_out <= r_48_27;
		if (write_en==1'b1)
			r_48_27 <= data_in;
	if (addr_selector[48]&addr_selector[28])
		data_out <= r_48_28;
		if (write_en==1'b1)
			r_48_28 <= data_in;
	if (addr_selector[48]&addr_selector[29])
		data_out <= r_48_29;
		if (write_en==1'b1)
			r_48_29 <= data_in;
	if (addr_selector[48]&addr_selector[30])
		data_out <= r_48_30;
		if (write_en==1'b1)
			r_48_30 <= data_in;
	if (addr_selector[48]&addr_selector[31])
		data_out <= r_48_31;
		if (write_en==1'b1)
			r_48_31 <= data_in;
	if (addr_selector[48]&addr_selector[32])
		data_out <= r_48_32;
		if (write_en==1'b1)
			r_48_32 <= data_in;
	if (addr_selector[48]&addr_selector[33])
		data_out <= r_48_33;
		if (write_en==1'b1)
			r_48_33 <= data_in;
	if (addr_selector[48]&addr_selector[34])
		data_out <= r_48_34;
		if (write_en==1'b1)
			r_48_34 <= data_in;
	if (addr_selector[48]&addr_selector[35])
		data_out <= r_48_35;
		if (write_en==1'b1)
			r_48_35 <= data_in;
	if (addr_selector[48]&addr_selector[36])
		data_out <= r_48_36;
		if (write_en==1'b1)
			r_48_36 <= data_in;
	if (addr_selector[48]&addr_selector[37])
		data_out <= r_48_37;
		if (write_en==1'b1)
			r_48_37 <= data_in;
	if (addr_selector[48]&addr_selector[38])
		data_out <= r_48_38;
		if (write_en==1'b1)
			r_48_38 <= data_in;
	if (addr_selector[48]&addr_selector[39])
		data_out <= r_48_39;
		if (write_en==1'b1)
			r_48_39 <= data_in;
	if (addr_selector[48]&addr_selector[40])
		data_out <= r_48_40;
		if (write_en==1'b1)
			r_48_40 <= data_in;
	if (addr_selector[48]&addr_selector[41])
		data_out <= r_48_41;
		if (write_en==1'b1)
			r_48_41 <= data_in;
	if (addr_selector[48]&addr_selector[42])
		data_out <= r_48_42;
		if (write_en==1'b1)
			r_48_42 <= data_in;
	if (addr_selector[48]&addr_selector[43])
		data_out <= r_48_43;
		if (write_en==1'b1)
			r_48_43 <= data_in;
	if (addr_selector[48]&addr_selector[44])
		data_out <= r_48_44;
		if (write_en==1'b1)
			r_48_44 <= data_in;
	if (addr_selector[48]&addr_selector[45])
		data_out <= r_48_45;
		if (write_en==1'b1)
			r_48_45 <= data_in;
	if (addr_selector[48]&addr_selector[46])
		data_out <= r_48_46;
		if (write_en==1'b1)
			r_48_46 <= data_in;
	if (addr_selector[48]&addr_selector[47])
		data_out <= r_48_47;
		if (write_en==1'b1)
			r_48_47 <= data_in;
	if (addr_selector[48]&addr_selector[48])
		data_out <= r_48_48;
		if (write_en==1'b1)
			r_48_48 <= data_in;
	if (addr_selector[48]&addr_selector[49])
		data_out <= r_48_49;
		if (write_en==1'b1)
			r_48_49 <= data_in;
	if (addr_selector[48]&addr_selector[50])
		data_out <= r_48_50;
		if (write_en==1'b1)
			r_48_50 <= data_in;
	if (addr_selector[48]&addr_selector[51])
		data_out <= r_48_51;
		if (write_en==1'b1)
			r_48_51 <= data_in;
	if (addr_selector[48]&addr_selector[52])
		data_out <= r_48_52;
		if (write_en==1'b1)
			r_48_52 <= data_in;
	if (addr_selector[48]&addr_selector[53])
		data_out <= r_48_53;
		if (write_en==1'b1)
			r_48_53 <= data_in;
	if (addr_selector[48]&addr_selector[54])
		data_out <= r_48_54;
		if (write_en==1'b1)
			r_48_54 <= data_in;
	if (addr_selector[48]&addr_selector[55])
		data_out <= r_48_55;
		if (write_en==1'b1)
			r_48_55 <= data_in;
	if (addr_selector[48]&addr_selector[56])
		data_out <= r_48_56;
		if (write_en==1'b1)
			r_48_56 <= data_in;
	if (addr_selector[48]&addr_selector[57])
		data_out <= r_48_57;
		if (write_en==1'b1)
			r_48_57 <= data_in;
	if (addr_selector[48]&addr_selector[58])
		data_out <= r_48_58;
		if (write_en==1'b1)
			r_48_58 <= data_in;
	if (addr_selector[48]&addr_selector[59])
		data_out <= r_48_59;
		if (write_en==1'b1)
			r_48_59 <= data_in;
	if (addr_selector[48]&addr_selector[60])
		data_out <= r_48_60;
		if (write_en==1'b1)
			r_48_60 <= data_in;
	if (addr_selector[48]&addr_selector[61])
		data_out <= r_48_61;
		if (write_en==1'b1)
			r_48_61 <= data_in;
	if (addr_selector[48]&addr_selector[62])
		data_out <= r_48_62;
		if (write_en==1'b1)
			r_48_62 <= data_in;
	if (addr_selector[48]&addr_selector[63])
		data_out <= r_48_63;
		if (write_en==1'b1)
			r_48_63 <= data_in;
	if (addr_selector[49]&addr_selector[0])
		data_out <= r_49_0;
		if (write_en==1'b1)
			r_49_0 <= data_in;
	if (addr_selector[49]&addr_selector[1])
		data_out <= r_49_1;
		if (write_en==1'b1)
			r_49_1 <= data_in;
	if (addr_selector[49]&addr_selector[2])
		data_out <= r_49_2;
		if (write_en==1'b1)
			r_49_2 <= data_in;
	if (addr_selector[49]&addr_selector[3])
		data_out <= r_49_3;
		if (write_en==1'b1)
			r_49_3 <= data_in;
	if (addr_selector[49]&addr_selector[4])
		data_out <= r_49_4;
		if (write_en==1'b1)
			r_49_4 <= data_in;
	if (addr_selector[49]&addr_selector[5])
		data_out <= r_49_5;
		if (write_en==1'b1)
			r_49_5 <= data_in;
	if (addr_selector[49]&addr_selector[6])
		data_out <= r_49_6;
		if (write_en==1'b1)
			r_49_6 <= data_in;
	if (addr_selector[49]&addr_selector[7])
		data_out <= r_49_7;
		if (write_en==1'b1)
			r_49_7 <= data_in;
	if (addr_selector[49]&addr_selector[8])
		data_out <= r_49_8;
		if (write_en==1'b1)
			r_49_8 <= data_in;
	if (addr_selector[49]&addr_selector[9])
		data_out <= r_49_9;
		if (write_en==1'b1)
			r_49_9 <= data_in;
	if (addr_selector[49]&addr_selector[10])
		data_out <= r_49_10;
		if (write_en==1'b1)
			r_49_10 <= data_in;
	if (addr_selector[49]&addr_selector[11])
		data_out <= r_49_11;
		if (write_en==1'b1)
			r_49_11 <= data_in;
	if (addr_selector[49]&addr_selector[12])
		data_out <= r_49_12;
		if (write_en==1'b1)
			r_49_12 <= data_in;
	if (addr_selector[49]&addr_selector[13])
		data_out <= r_49_13;
		if (write_en==1'b1)
			r_49_13 <= data_in;
	if (addr_selector[49]&addr_selector[14])
		data_out <= r_49_14;
		if (write_en==1'b1)
			r_49_14 <= data_in;
	if (addr_selector[49]&addr_selector[15])
		data_out <= r_49_15;
		if (write_en==1'b1)
			r_49_15 <= data_in;
	if (addr_selector[49]&addr_selector[16])
		data_out <= r_49_16;
		if (write_en==1'b1)
			r_49_16 <= data_in;
	if (addr_selector[49]&addr_selector[17])
		data_out <= r_49_17;
		if (write_en==1'b1)
			r_49_17 <= data_in;
	if (addr_selector[49]&addr_selector[18])
		data_out <= r_49_18;
		if (write_en==1'b1)
			r_49_18 <= data_in;
	if (addr_selector[49]&addr_selector[19])
		data_out <= r_49_19;
		if (write_en==1'b1)
			r_49_19 <= data_in;
	if (addr_selector[49]&addr_selector[20])
		data_out <= r_49_20;
		if (write_en==1'b1)
			r_49_20 <= data_in;
	if (addr_selector[49]&addr_selector[21])
		data_out <= r_49_21;
		if (write_en==1'b1)
			r_49_21 <= data_in;
	if (addr_selector[49]&addr_selector[22])
		data_out <= r_49_22;
		if (write_en==1'b1)
			r_49_22 <= data_in;
	if (addr_selector[49]&addr_selector[23])
		data_out <= r_49_23;
		if (write_en==1'b1)
			r_49_23 <= data_in;
	if (addr_selector[49]&addr_selector[24])
		data_out <= r_49_24;
		if (write_en==1'b1)
			r_49_24 <= data_in;
	if (addr_selector[49]&addr_selector[25])
		data_out <= r_49_25;
		if (write_en==1'b1)
			r_49_25 <= data_in;
	if (addr_selector[49]&addr_selector[26])
		data_out <= r_49_26;
		if (write_en==1'b1)
			r_49_26 <= data_in;
	if (addr_selector[49]&addr_selector[27])
		data_out <= r_49_27;
		if (write_en==1'b1)
			r_49_27 <= data_in;
	if (addr_selector[49]&addr_selector[28])
		data_out <= r_49_28;
		if (write_en==1'b1)
			r_49_28 <= data_in;
	if (addr_selector[49]&addr_selector[29])
		data_out <= r_49_29;
		if (write_en==1'b1)
			r_49_29 <= data_in;
	if (addr_selector[49]&addr_selector[30])
		data_out <= r_49_30;
		if (write_en==1'b1)
			r_49_30 <= data_in;
	if (addr_selector[49]&addr_selector[31])
		data_out <= r_49_31;
		if (write_en==1'b1)
			r_49_31 <= data_in;
	if (addr_selector[49]&addr_selector[32])
		data_out <= r_49_32;
		if (write_en==1'b1)
			r_49_32 <= data_in;
	if (addr_selector[49]&addr_selector[33])
		data_out <= r_49_33;
		if (write_en==1'b1)
			r_49_33 <= data_in;
	if (addr_selector[49]&addr_selector[34])
		data_out <= r_49_34;
		if (write_en==1'b1)
			r_49_34 <= data_in;
	if (addr_selector[49]&addr_selector[35])
		data_out <= r_49_35;
		if (write_en==1'b1)
			r_49_35 <= data_in;
	if (addr_selector[49]&addr_selector[36])
		data_out <= r_49_36;
		if (write_en==1'b1)
			r_49_36 <= data_in;
	if (addr_selector[49]&addr_selector[37])
		data_out <= r_49_37;
		if (write_en==1'b1)
			r_49_37 <= data_in;
	if (addr_selector[49]&addr_selector[38])
		data_out <= r_49_38;
		if (write_en==1'b1)
			r_49_38 <= data_in;
	if (addr_selector[49]&addr_selector[39])
		data_out <= r_49_39;
		if (write_en==1'b1)
			r_49_39 <= data_in;
	if (addr_selector[49]&addr_selector[40])
		data_out <= r_49_40;
		if (write_en==1'b1)
			r_49_40 <= data_in;
	if (addr_selector[49]&addr_selector[41])
		data_out <= r_49_41;
		if (write_en==1'b1)
			r_49_41 <= data_in;
	if (addr_selector[49]&addr_selector[42])
		data_out <= r_49_42;
		if (write_en==1'b1)
			r_49_42 <= data_in;
	if (addr_selector[49]&addr_selector[43])
		data_out <= r_49_43;
		if (write_en==1'b1)
			r_49_43 <= data_in;
	if (addr_selector[49]&addr_selector[44])
		data_out <= r_49_44;
		if (write_en==1'b1)
			r_49_44 <= data_in;
	if (addr_selector[49]&addr_selector[45])
		data_out <= r_49_45;
		if (write_en==1'b1)
			r_49_45 <= data_in;
	if (addr_selector[49]&addr_selector[46])
		data_out <= r_49_46;
		if (write_en==1'b1)
			r_49_46 <= data_in;
	if (addr_selector[49]&addr_selector[47])
		data_out <= r_49_47;
		if (write_en==1'b1)
			r_49_47 <= data_in;
	if (addr_selector[49]&addr_selector[48])
		data_out <= r_49_48;
		if (write_en==1'b1)
			r_49_48 <= data_in;
	if (addr_selector[49]&addr_selector[49])
		data_out <= r_49_49;
		if (write_en==1'b1)
			r_49_49 <= data_in;
	if (addr_selector[49]&addr_selector[50])
		data_out <= r_49_50;
		if (write_en==1'b1)
			r_49_50 <= data_in;
	if (addr_selector[49]&addr_selector[51])
		data_out <= r_49_51;
		if (write_en==1'b1)
			r_49_51 <= data_in;
	if (addr_selector[49]&addr_selector[52])
		data_out <= r_49_52;
		if (write_en==1'b1)
			r_49_52 <= data_in;
	if (addr_selector[49]&addr_selector[53])
		data_out <= r_49_53;
		if (write_en==1'b1)
			r_49_53 <= data_in;
	if (addr_selector[49]&addr_selector[54])
		data_out <= r_49_54;
		if (write_en==1'b1)
			r_49_54 <= data_in;
	if (addr_selector[49]&addr_selector[55])
		data_out <= r_49_55;
		if (write_en==1'b1)
			r_49_55 <= data_in;
	if (addr_selector[49]&addr_selector[56])
		data_out <= r_49_56;
		if (write_en==1'b1)
			r_49_56 <= data_in;
	if (addr_selector[49]&addr_selector[57])
		data_out <= r_49_57;
		if (write_en==1'b1)
			r_49_57 <= data_in;
	if (addr_selector[49]&addr_selector[58])
		data_out <= r_49_58;
		if (write_en==1'b1)
			r_49_58 <= data_in;
	if (addr_selector[49]&addr_selector[59])
		data_out <= r_49_59;
		if (write_en==1'b1)
			r_49_59 <= data_in;
	if (addr_selector[49]&addr_selector[60])
		data_out <= r_49_60;
		if (write_en==1'b1)
			r_49_60 <= data_in;
	if (addr_selector[49]&addr_selector[61])
		data_out <= r_49_61;
		if (write_en==1'b1)
			r_49_61 <= data_in;
	if (addr_selector[49]&addr_selector[62])
		data_out <= r_49_62;
		if (write_en==1'b1)
			r_49_62 <= data_in;
	if (addr_selector[49]&addr_selector[63])
		data_out <= r_49_63;
		if (write_en==1'b1)
			r_49_63 <= data_in;
	if (addr_selector[50]&addr_selector[0])
		data_out <= r_50_0;
		if (write_en==1'b1)
			r_50_0 <= data_in;
	if (addr_selector[50]&addr_selector[1])
		data_out <= r_50_1;
		if (write_en==1'b1)
			r_50_1 <= data_in;
	if (addr_selector[50]&addr_selector[2])
		data_out <= r_50_2;
		if (write_en==1'b1)
			r_50_2 <= data_in;
	if (addr_selector[50]&addr_selector[3])
		data_out <= r_50_3;
		if (write_en==1'b1)
			r_50_3 <= data_in;
	if (addr_selector[50]&addr_selector[4])
		data_out <= r_50_4;
		if (write_en==1'b1)
			r_50_4 <= data_in;
	if (addr_selector[50]&addr_selector[5])
		data_out <= r_50_5;
		if (write_en==1'b1)
			r_50_5 <= data_in;
	if (addr_selector[50]&addr_selector[6])
		data_out <= r_50_6;
		if (write_en==1'b1)
			r_50_6 <= data_in;
	if (addr_selector[50]&addr_selector[7])
		data_out <= r_50_7;
		if (write_en==1'b1)
			r_50_7 <= data_in;
	if (addr_selector[50]&addr_selector[8])
		data_out <= r_50_8;
		if (write_en==1'b1)
			r_50_8 <= data_in;
	if (addr_selector[50]&addr_selector[9])
		data_out <= r_50_9;
		if (write_en==1'b1)
			r_50_9 <= data_in;
	if (addr_selector[50]&addr_selector[10])
		data_out <= r_50_10;
		if (write_en==1'b1)
			r_50_10 <= data_in;
	if (addr_selector[50]&addr_selector[11])
		data_out <= r_50_11;
		if (write_en==1'b1)
			r_50_11 <= data_in;
	if (addr_selector[50]&addr_selector[12])
		data_out <= r_50_12;
		if (write_en==1'b1)
			r_50_12 <= data_in;
	if (addr_selector[50]&addr_selector[13])
		data_out <= r_50_13;
		if (write_en==1'b1)
			r_50_13 <= data_in;
	if (addr_selector[50]&addr_selector[14])
		data_out <= r_50_14;
		if (write_en==1'b1)
			r_50_14 <= data_in;
	if (addr_selector[50]&addr_selector[15])
		data_out <= r_50_15;
		if (write_en==1'b1)
			r_50_15 <= data_in;
	if (addr_selector[50]&addr_selector[16])
		data_out <= r_50_16;
		if (write_en==1'b1)
			r_50_16 <= data_in;
	if (addr_selector[50]&addr_selector[17])
		data_out <= r_50_17;
		if (write_en==1'b1)
			r_50_17 <= data_in;
	if (addr_selector[50]&addr_selector[18])
		data_out <= r_50_18;
		if (write_en==1'b1)
			r_50_18 <= data_in;
	if (addr_selector[50]&addr_selector[19])
		data_out <= r_50_19;
		if (write_en==1'b1)
			r_50_19 <= data_in;
	if (addr_selector[50]&addr_selector[20])
		data_out <= r_50_20;
		if (write_en==1'b1)
			r_50_20 <= data_in;
	if (addr_selector[50]&addr_selector[21])
		data_out <= r_50_21;
		if (write_en==1'b1)
			r_50_21 <= data_in;
	if (addr_selector[50]&addr_selector[22])
		data_out <= r_50_22;
		if (write_en==1'b1)
			r_50_22 <= data_in;
	if (addr_selector[50]&addr_selector[23])
		data_out <= r_50_23;
		if (write_en==1'b1)
			r_50_23 <= data_in;
	if (addr_selector[50]&addr_selector[24])
		data_out <= r_50_24;
		if (write_en==1'b1)
			r_50_24 <= data_in;
	if (addr_selector[50]&addr_selector[25])
		data_out <= r_50_25;
		if (write_en==1'b1)
			r_50_25 <= data_in;
	if (addr_selector[50]&addr_selector[26])
		data_out <= r_50_26;
		if (write_en==1'b1)
			r_50_26 <= data_in;
	if (addr_selector[50]&addr_selector[27])
		data_out <= r_50_27;
		if (write_en==1'b1)
			r_50_27 <= data_in;
	if (addr_selector[50]&addr_selector[28])
		data_out <= r_50_28;
		if (write_en==1'b1)
			r_50_28 <= data_in;
	if (addr_selector[50]&addr_selector[29])
		data_out <= r_50_29;
		if (write_en==1'b1)
			r_50_29 <= data_in;
	if (addr_selector[50]&addr_selector[30])
		data_out <= r_50_30;
		if (write_en==1'b1)
			r_50_30 <= data_in;
	if (addr_selector[50]&addr_selector[31])
		data_out <= r_50_31;
		if (write_en==1'b1)
			r_50_31 <= data_in;
	if (addr_selector[50]&addr_selector[32])
		data_out <= r_50_32;
		if (write_en==1'b1)
			r_50_32 <= data_in;
	if (addr_selector[50]&addr_selector[33])
		data_out <= r_50_33;
		if (write_en==1'b1)
			r_50_33 <= data_in;
	if (addr_selector[50]&addr_selector[34])
		data_out <= r_50_34;
		if (write_en==1'b1)
			r_50_34 <= data_in;
	if (addr_selector[50]&addr_selector[35])
		data_out <= r_50_35;
		if (write_en==1'b1)
			r_50_35 <= data_in;
	if (addr_selector[50]&addr_selector[36])
		data_out <= r_50_36;
		if (write_en==1'b1)
			r_50_36 <= data_in;
	if (addr_selector[50]&addr_selector[37])
		data_out <= r_50_37;
		if (write_en==1'b1)
			r_50_37 <= data_in;
	if (addr_selector[50]&addr_selector[38])
		data_out <= r_50_38;
		if (write_en==1'b1)
			r_50_38 <= data_in;
	if (addr_selector[50]&addr_selector[39])
		data_out <= r_50_39;
		if (write_en==1'b1)
			r_50_39 <= data_in;
	if (addr_selector[50]&addr_selector[40])
		data_out <= r_50_40;
		if (write_en==1'b1)
			r_50_40 <= data_in;
	if (addr_selector[50]&addr_selector[41])
		data_out <= r_50_41;
		if (write_en==1'b1)
			r_50_41 <= data_in;
	if (addr_selector[50]&addr_selector[42])
		data_out <= r_50_42;
		if (write_en==1'b1)
			r_50_42 <= data_in;
	if (addr_selector[50]&addr_selector[43])
		data_out <= r_50_43;
		if (write_en==1'b1)
			r_50_43 <= data_in;
	if (addr_selector[50]&addr_selector[44])
		data_out <= r_50_44;
		if (write_en==1'b1)
			r_50_44 <= data_in;
	if (addr_selector[50]&addr_selector[45])
		data_out <= r_50_45;
		if (write_en==1'b1)
			r_50_45 <= data_in;
	if (addr_selector[50]&addr_selector[46])
		data_out <= r_50_46;
		if (write_en==1'b1)
			r_50_46 <= data_in;
	if (addr_selector[50]&addr_selector[47])
		data_out <= r_50_47;
		if (write_en==1'b1)
			r_50_47 <= data_in;
	if (addr_selector[50]&addr_selector[48])
		data_out <= r_50_48;
		if (write_en==1'b1)
			r_50_48 <= data_in;
	if (addr_selector[50]&addr_selector[49])
		data_out <= r_50_49;
		if (write_en==1'b1)
			r_50_49 <= data_in;
	if (addr_selector[50]&addr_selector[50])
		data_out <= r_50_50;
		if (write_en==1'b1)
			r_50_50 <= data_in;
	if (addr_selector[50]&addr_selector[51])
		data_out <= r_50_51;
		if (write_en==1'b1)
			r_50_51 <= data_in;
	if (addr_selector[50]&addr_selector[52])
		data_out <= r_50_52;
		if (write_en==1'b1)
			r_50_52 <= data_in;
	if (addr_selector[50]&addr_selector[53])
		data_out <= r_50_53;
		if (write_en==1'b1)
			r_50_53 <= data_in;
	if (addr_selector[50]&addr_selector[54])
		data_out <= r_50_54;
		if (write_en==1'b1)
			r_50_54 <= data_in;
	if (addr_selector[50]&addr_selector[55])
		data_out <= r_50_55;
		if (write_en==1'b1)
			r_50_55 <= data_in;
	if (addr_selector[50]&addr_selector[56])
		data_out <= r_50_56;
		if (write_en==1'b1)
			r_50_56 <= data_in;
	if (addr_selector[50]&addr_selector[57])
		data_out <= r_50_57;
		if (write_en==1'b1)
			r_50_57 <= data_in;
	if (addr_selector[50]&addr_selector[58])
		data_out <= r_50_58;
		if (write_en==1'b1)
			r_50_58 <= data_in;
	if (addr_selector[50]&addr_selector[59])
		data_out <= r_50_59;
		if (write_en==1'b1)
			r_50_59 <= data_in;
	if (addr_selector[50]&addr_selector[60])
		data_out <= r_50_60;
		if (write_en==1'b1)
			r_50_60 <= data_in;
	if (addr_selector[50]&addr_selector[61])
		data_out <= r_50_61;
		if (write_en==1'b1)
			r_50_61 <= data_in;
	if (addr_selector[50]&addr_selector[62])
		data_out <= r_50_62;
		if (write_en==1'b1)
			r_50_62 <= data_in;
	if (addr_selector[50]&addr_selector[63])
		data_out <= r_50_63;
		if (write_en==1'b1)
			r_50_63 <= data_in;
	if (addr_selector[51]&addr_selector[0])
		data_out <= r_51_0;
		if (write_en==1'b1)
			r_51_0 <= data_in;
	if (addr_selector[51]&addr_selector[1])
		data_out <= r_51_1;
		if (write_en==1'b1)
			r_51_1 <= data_in;
	if (addr_selector[51]&addr_selector[2])
		data_out <= r_51_2;
		if (write_en==1'b1)
			r_51_2 <= data_in;
	if (addr_selector[51]&addr_selector[3])
		data_out <= r_51_3;
		if (write_en==1'b1)
			r_51_3 <= data_in;
	if (addr_selector[51]&addr_selector[4])
		data_out <= r_51_4;
		if (write_en==1'b1)
			r_51_4 <= data_in;
	if (addr_selector[51]&addr_selector[5])
		data_out <= r_51_5;
		if (write_en==1'b1)
			r_51_5 <= data_in;
	if (addr_selector[51]&addr_selector[6])
		data_out <= r_51_6;
		if (write_en==1'b1)
			r_51_6 <= data_in;
	if (addr_selector[51]&addr_selector[7])
		data_out <= r_51_7;
		if (write_en==1'b1)
			r_51_7 <= data_in;
	if (addr_selector[51]&addr_selector[8])
		data_out <= r_51_8;
		if (write_en==1'b1)
			r_51_8 <= data_in;
	if (addr_selector[51]&addr_selector[9])
		data_out <= r_51_9;
		if (write_en==1'b1)
			r_51_9 <= data_in;
	if (addr_selector[51]&addr_selector[10])
		data_out <= r_51_10;
		if (write_en==1'b1)
			r_51_10 <= data_in;
	if (addr_selector[51]&addr_selector[11])
		data_out <= r_51_11;
		if (write_en==1'b1)
			r_51_11 <= data_in;
	if (addr_selector[51]&addr_selector[12])
		data_out <= r_51_12;
		if (write_en==1'b1)
			r_51_12 <= data_in;
	if (addr_selector[51]&addr_selector[13])
		data_out <= r_51_13;
		if (write_en==1'b1)
			r_51_13 <= data_in;
	if (addr_selector[51]&addr_selector[14])
		data_out <= r_51_14;
		if (write_en==1'b1)
			r_51_14 <= data_in;
	if (addr_selector[51]&addr_selector[15])
		data_out <= r_51_15;
		if (write_en==1'b1)
			r_51_15 <= data_in;
	if (addr_selector[51]&addr_selector[16])
		data_out <= r_51_16;
		if (write_en==1'b1)
			r_51_16 <= data_in;
	if (addr_selector[51]&addr_selector[17])
		data_out <= r_51_17;
		if (write_en==1'b1)
			r_51_17 <= data_in;
	if (addr_selector[51]&addr_selector[18])
		data_out <= r_51_18;
		if (write_en==1'b1)
			r_51_18 <= data_in;
	if (addr_selector[51]&addr_selector[19])
		data_out <= r_51_19;
		if (write_en==1'b1)
			r_51_19 <= data_in;
	if (addr_selector[51]&addr_selector[20])
		data_out <= r_51_20;
		if (write_en==1'b1)
			r_51_20 <= data_in;
	if (addr_selector[51]&addr_selector[21])
		data_out <= r_51_21;
		if (write_en==1'b1)
			r_51_21 <= data_in;
	if (addr_selector[51]&addr_selector[22])
		data_out <= r_51_22;
		if (write_en==1'b1)
			r_51_22 <= data_in;
	if (addr_selector[51]&addr_selector[23])
		data_out <= r_51_23;
		if (write_en==1'b1)
			r_51_23 <= data_in;
	if (addr_selector[51]&addr_selector[24])
		data_out <= r_51_24;
		if (write_en==1'b1)
			r_51_24 <= data_in;
	if (addr_selector[51]&addr_selector[25])
		data_out <= r_51_25;
		if (write_en==1'b1)
			r_51_25 <= data_in;
	if (addr_selector[51]&addr_selector[26])
		data_out <= r_51_26;
		if (write_en==1'b1)
			r_51_26 <= data_in;
	if (addr_selector[51]&addr_selector[27])
		data_out <= r_51_27;
		if (write_en==1'b1)
			r_51_27 <= data_in;
	if (addr_selector[51]&addr_selector[28])
		data_out <= r_51_28;
		if (write_en==1'b1)
			r_51_28 <= data_in;
	if (addr_selector[51]&addr_selector[29])
		data_out <= r_51_29;
		if (write_en==1'b1)
			r_51_29 <= data_in;
	if (addr_selector[51]&addr_selector[30])
		data_out <= r_51_30;
		if (write_en==1'b1)
			r_51_30 <= data_in;
	if (addr_selector[51]&addr_selector[31])
		data_out <= r_51_31;
		if (write_en==1'b1)
			r_51_31 <= data_in;
	if (addr_selector[51]&addr_selector[32])
		data_out <= r_51_32;
		if (write_en==1'b1)
			r_51_32 <= data_in;
	if (addr_selector[51]&addr_selector[33])
		data_out <= r_51_33;
		if (write_en==1'b1)
			r_51_33 <= data_in;
	if (addr_selector[51]&addr_selector[34])
		data_out <= r_51_34;
		if (write_en==1'b1)
			r_51_34 <= data_in;
	if (addr_selector[51]&addr_selector[35])
		data_out <= r_51_35;
		if (write_en==1'b1)
			r_51_35 <= data_in;
	if (addr_selector[51]&addr_selector[36])
		data_out <= r_51_36;
		if (write_en==1'b1)
			r_51_36 <= data_in;
	if (addr_selector[51]&addr_selector[37])
		data_out <= r_51_37;
		if (write_en==1'b1)
			r_51_37 <= data_in;
	if (addr_selector[51]&addr_selector[38])
		data_out <= r_51_38;
		if (write_en==1'b1)
			r_51_38 <= data_in;
	if (addr_selector[51]&addr_selector[39])
		data_out <= r_51_39;
		if (write_en==1'b1)
			r_51_39 <= data_in;
	if (addr_selector[51]&addr_selector[40])
		data_out <= r_51_40;
		if (write_en==1'b1)
			r_51_40 <= data_in;
	if (addr_selector[51]&addr_selector[41])
		data_out <= r_51_41;
		if (write_en==1'b1)
			r_51_41 <= data_in;
	if (addr_selector[51]&addr_selector[42])
		data_out <= r_51_42;
		if (write_en==1'b1)
			r_51_42 <= data_in;
	if (addr_selector[51]&addr_selector[43])
		data_out <= r_51_43;
		if (write_en==1'b1)
			r_51_43 <= data_in;
	if (addr_selector[51]&addr_selector[44])
		data_out <= r_51_44;
		if (write_en==1'b1)
			r_51_44 <= data_in;
	if (addr_selector[51]&addr_selector[45])
		data_out <= r_51_45;
		if (write_en==1'b1)
			r_51_45 <= data_in;
	if (addr_selector[51]&addr_selector[46])
		data_out <= r_51_46;
		if (write_en==1'b1)
			r_51_46 <= data_in;
	if (addr_selector[51]&addr_selector[47])
		data_out <= r_51_47;
		if (write_en==1'b1)
			r_51_47 <= data_in;
	if (addr_selector[51]&addr_selector[48])
		data_out <= r_51_48;
		if (write_en==1'b1)
			r_51_48 <= data_in;
	if (addr_selector[51]&addr_selector[49])
		data_out <= r_51_49;
		if (write_en==1'b1)
			r_51_49 <= data_in;
	if (addr_selector[51]&addr_selector[50])
		data_out <= r_51_50;
		if (write_en==1'b1)
			r_51_50 <= data_in;
	if (addr_selector[51]&addr_selector[51])
		data_out <= r_51_51;
		if (write_en==1'b1)
			r_51_51 <= data_in;
	if (addr_selector[51]&addr_selector[52])
		data_out <= r_51_52;
		if (write_en==1'b1)
			r_51_52 <= data_in;
	if (addr_selector[51]&addr_selector[53])
		data_out <= r_51_53;
		if (write_en==1'b1)
			r_51_53 <= data_in;
	if (addr_selector[51]&addr_selector[54])
		data_out <= r_51_54;
		if (write_en==1'b1)
			r_51_54 <= data_in;
	if (addr_selector[51]&addr_selector[55])
		data_out <= r_51_55;
		if (write_en==1'b1)
			r_51_55 <= data_in;
	if (addr_selector[51]&addr_selector[56])
		data_out <= r_51_56;
		if (write_en==1'b1)
			r_51_56 <= data_in;
	if (addr_selector[51]&addr_selector[57])
		data_out <= r_51_57;
		if (write_en==1'b1)
			r_51_57 <= data_in;
	if (addr_selector[51]&addr_selector[58])
		data_out <= r_51_58;
		if (write_en==1'b1)
			r_51_58 <= data_in;
	if (addr_selector[51]&addr_selector[59])
		data_out <= r_51_59;
		if (write_en==1'b1)
			r_51_59 <= data_in;
	if (addr_selector[51]&addr_selector[60])
		data_out <= r_51_60;
		if (write_en==1'b1)
			r_51_60 <= data_in;
	if (addr_selector[51]&addr_selector[61])
		data_out <= r_51_61;
		if (write_en==1'b1)
			r_51_61 <= data_in;
	if (addr_selector[51]&addr_selector[62])
		data_out <= r_51_62;
		if (write_en==1'b1)
			r_51_62 <= data_in;
	if (addr_selector[51]&addr_selector[63])
		data_out <= r_51_63;
		if (write_en==1'b1)
			r_51_63 <= data_in;
	if (addr_selector[52]&addr_selector[0])
		data_out <= r_52_0;
		if (write_en==1'b1)
			r_52_0 <= data_in;
	if (addr_selector[52]&addr_selector[1])
		data_out <= r_52_1;
		if (write_en==1'b1)
			r_52_1 <= data_in;
	if (addr_selector[52]&addr_selector[2])
		data_out <= r_52_2;
		if (write_en==1'b1)
			r_52_2 <= data_in;
	if (addr_selector[52]&addr_selector[3])
		data_out <= r_52_3;
		if (write_en==1'b1)
			r_52_3 <= data_in;
	if (addr_selector[52]&addr_selector[4])
		data_out <= r_52_4;
		if (write_en==1'b1)
			r_52_4 <= data_in;
	if (addr_selector[52]&addr_selector[5])
		data_out <= r_52_5;
		if (write_en==1'b1)
			r_52_5 <= data_in;
	if (addr_selector[52]&addr_selector[6])
		data_out <= r_52_6;
		if (write_en==1'b1)
			r_52_6 <= data_in;
	if (addr_selector[52]&addr_selector[7])
		data_out <= r_52_7;
		if (write_en==1'b1)
			r_52_7 <= data_in;
	if (addr_selector[52]&addr_selector[8])
		data_out <= r_52_8;
		if (write_en==1'b1)
			r_52_8 <= data_in;
	if (addr_selector[52]&addr_selector[9])
		data_out <= r_52_9;
		if (write_en==1'b1)
			r_52_9 <= data_in;
	if (addr_selector[52]&addr_selector[10])
		data_out <= r_52_10;
		if (write_en==1'b1)
			r_52_10 <= data_in;
	if (addr_selector[52]&addr_selector[11])
		data_out <= r_52_11;
		if (write_en==1'b1)
			r_52_11 <= data_in;
	if (addr_selector[52]&addr_selector[12])
		data_out <= r_52_12;
		if (write_en==1'b1)
			r_52_12 <= data_in;
	if (addr_selector[52]&addr_selector[13])
		data_out <= r_52_13;
		if (write_en==1'b1)
			r_52_13 <= data_in;
	if (addr_selector[52]&addr_selector[14])
		data_out <= r_52_14;
		if (write_en==1'b1)
			r_52_14 <= data_in;
	if (addr_selector[52]&addr_selector[15])
		data_out <= r_52_15;
		if (write_en==1'b1)
			r_52_15 <= data_in;
	if (addr_selector[52]&addr_selector[16])
		data_out <= r_52_16;
		if (write_en==1'b1)
			r_52_16 <= data_in;
	if (addr_selector[52]&addr_selector[17])
		data_out <= r_52_17;
		if (write_en==1'b1)
			r_52_17 <= data_in;
	if (addr_selector[52]&addr_selector[18])
		data_out <= r_52_18;
		if (write_en==1'b1)
			r_52_18 <= data_in;
	if (addr_selector[52]&addr_selector[19])
		data_out <= r_52_19;
		if (write_en==1'b1)
			r_52_19 <= data_in;
	if (addr_selector[52]&addr_selector[20])
		data_out <= r_52_20;
		if (write_en==1'b1)
			r_52_20 <= data_in;
	if (addr_selector[52]&addr_selector[21])
		data_out <= r_52_21;
		if (write_en==1'b1)
			r_52_21 <= data_in;
	if (addr_selector[52]&addr_selector[22])
		data_out <= r_52_22;
		if (write_en==1'b1)
			r_52_22 <= data_in;
	if (addr_selector[52]&addr_selector[23])
		data_out <= r_52_23;
		if (write_en==1'b1)
			r_52_23 <= data_in;
	if (addr_selector[52]&addr_selector[24])
		data_out <= r_52_24;
		if (write_en==1'b1)
			r_52_24 <= data_in;
	if (addr_selector[52]&addr_selector[25])
		data_out <= r_52_25;
		if (write_en==1'b1)
			r_52_25 <= data_in;
	if (addr_selector[52]&addr_selector[26])
		data_out <= r_52_26;
		if (write_en==1'b1)
			r_52_26 <= data_in;
	if (addr_selector[52]&addr_selector[27])
		data_out <= r_52_27;
		if (write_en==1'b1)
			r_52_27 <= data_in;
	if (addr_selector[52]&addr_selector[28])
		data_out <= r_52_28;
		if (write_en==1'b1)
			r_52_28 <= data_in;
	if (addr_selector[52]&addr_selector[29])
		data_out <= r_52_29;
		if (write_en==1'b1)
			r_52_29 <= data_in;
	if (addr_selector[52]&addr_selector[30])
		data_out <= r_52_30;
		if (write_en==1'b1)
			r_52_30 <= data_in;
	if (addr_selector[52]&addr_selector[31])
		data_out <= r_52_31;
		if (write_en==1'b1)
			r_52_31 <= data_in;
	if (addr_selector[52]&addr_selector[32])
		data_out <= r_52_32;
		if (write_en==1'b1)
			r_52_32 <= data_in;
	if (addr_selector[52]&addr_selector[33])
		data_out <= r_52_33;
		if (write_en==1'b1)
			r_52_33 <= data_in;
	if (addr_selector[52]&addr_selector[34])
		data_out <= r_52_34;
		if (write_en==1'b1)
			r_52_34 <= data_in;
	if (addr_selector[52]&addr_selector[35])
		data_out <= r_52_35;
		if (write_en==1'b1)
			r_52_35 <= data_in;
	if (addr_selector[52]&addr_selector[36])
		data_out <= r_52_36;
		if (write_en==1'b1)
			r_52_36 <= data_in;
	if (addr_selector[52]&addr_selector[37])
		data_out <= r_52_37;
		if (write_en==1'b1)
			r_52_37 <= data_in;
	if (addr_selector[52]&addr_selector[38])
		data_out <= r_52_38;
		if (write_en==1'b1)
			r_52_38 <= data_in;
	if (addr_selector[52]&addr_selector[39])
		data_out <= r_52_39;
		if (write_en==1'b1)
			r_52_39 <= data_in;
	if (addr_selector[52]&addr_selector[40])
		data_out <= r_52_40;
		if (write_en==1'b1)
			r_52_40 <= data_in;
	if (addr_selector[52]&addr_selector[41])
		data_out <= r_52_41;
		if (write_en==1'b1)
			r_52_41 <= data_in;
	if (addr_selector[52]&addr_selector[42])
		data_out <= r_52_42;
		if (write_en==1'b1)
			r_52_42 <= data_in;
	if (addr_selector[52]&addr_selector[43])
		data_out <= r_52_43;
		if (write_en==1'b1)
			r_52_43 <= data_in;
	if (addr_selector[52]&addr_selector[44])
		data_out <= r_52_44;
		if (write_en==1'b1)
			r_52_44 <= data_in;
	if (addr_selector[52]&addr_selector[45])
		data_out <= r_52_45;
		if (write_en==1'b1)
			r_52_45 <= data_in;
	if (addr_selector[52]&addr_selector[46])
		data_out <= r_52_46;
		if (write_en==1'b1)
			r_52_46 <= data_in;
	if (addr_selector[52]&addr_selector[47])
		data_out <= r_52_47;
		if (write_en==1'b1)
			r_52_47 <= data_in;
	if (addr_selector[52]&addr_selector[48])
		data_out <= r_52_48;
		if (write_en==1'b1)
			r_52_48 <= data_in;
	if (addr_selector[52]&addr_selector[49])
		data_out <= r_52_49;
		if (write_en==1'b1)
			r_52_49 <= data_in;
	if (addr_selector[52]&addr_selector[50])
		data_out <= r_52_50;
		if (write_en==1'b1)
			r_52_50 <= data_in;
	if (addr_selector[52]&addr_selector[51])
		data_out <= r_52_51;
		if (write_en==1'b1)
			r_52_51 <= data_in;
	if (addr_selector[52]&addr_selector[52])
		data_out <= r_52_52;
		if (write_en==1'b1)
			r_52_52 <= data_in;
	if (addr_selector[52]&addr_selector[53])
		data_out <= r_52_53;
		if (write_en==1'b1)
			r_52_53 <= data_in;
	if (addr_selector[52]&addr_selector[54])
		data_out <= r_52_54;
		if (write_en==1'b1)
			r_52_54 <= data_in;
	if (addr_selector[52]&addr_selector[55])
		data_out <= r_52_55;
		if (write_en==1'b1)
			r_52_55 <= data_in;
	if (addr_selector[52]&addr_selector[56])
		data_out <= r_52_56;
		if (write_en==1'b1)
			r_52_56 <= data_in;
	if (addr_selector[52]&addr_selector[57])
		data_out <= r_52_57;
		if (write_en==1'b1)
			r_52_57 <= data_in;
	if (addr_selector[52]&addr_selector[58])
		data_out <= r_52_58;
		if (write_en==1'b1)
			r_52_58 <= data_in;
	if (addr_selector[52]&addr_selector[59])
		data_out <= r_52_59;
		if (write_en==1'b1)
			r_52_59 <= data_in;
	if (addr_selector[52]&addr_selector[60])
		data_out <= r_52_60;
		if (write_en==1'b1)
			r_52_60 <= data_in;
	if (addr_selector[52]&addr_selector[61])
		data_out <= r_52_61;
		if (write_en==1'b1)
			r_52_61 <= data_in;
	if (addr_selector[52]&addr_selector[62])
		data_out <= r_52_62;
		if (write_en==1'b1)
			r_52_62 <= data_in;
	if (addr_selector[52]&addr_selector[63])
		data_out <= r_52_63;
		if (write_en==1'b1)
			r_52_63 <= data_in;
	if (addr_selector[53]&addr_selector[0])
		data_out <= r_53_0;
		if (write_en==1'b1)
			r_53_0 <= data_in;
	if (addr_selector[53]&addr_selector[1])
		data_out <= r_53_1;
		if (write_en==1'b1)
			r_53_1 <= data_in;
	if (addr_selector[53]&addr_selector[2])
		data_out <= r_53_2;
		if (write_en==1'b1)
			r_53_2 <= data_in;
	if (addr_selector[53]&addr_selector[3])
		data_out <= r_53_3;
		if (write_en==1'b1)
			r_53_3 <= data_in;
	if (addr_selector[53]&addr_selector[4])
		data_out <= r_53_4;
		if (write_en==1'b1)
			r_53_4 <= data_in;
	if (addr_selector[53]&addr_selector[5])
		data_out <= r_53_5;
		if (write_en==1'b1)
			r_53_5 <= data_in;
	if (addr_selector[53]&addr_selector[6])
		data_out <= r_53_6;
		if (write_en==1'b1)
			r_53_6 <= data_in;
	if (addr_selector[53]&addr_selector[7])
		data_out <= r_53_7;
		if (write_en==1'b1)
			r_53_7 <= data_in;
	if (addr_selector[53]&addr_selector[8])
		data_out <= r_53_8;
		if (write_en==1'b1)
			r_53_8 <= data_in;
	if (addr_selector[53]&addr_selector[9])
		data_out <= r_53_9;
		if (write_en==1'b1)
			r_53_9 <= data_in;
	if (addr_selector[53]&addr_selector[10])
		data_out <= r_53_10;
		if (write_en==1'b1)
			r_53_10 <= data_in;
	if (addr_selector[53]&addr_selector[11])
		data_out <= r_53_11;
		if (write_en==1'b1)
			r_53_11 <= data_in;
	if (addr_selector[53]&addr_selector[12])
		data_out <= r_53_12;
		if (write_en==1'b1)
			r_53_12 <= data_in;
	if (addr_selector[53]&addr_selector[13])
		data_out <= r_53_13;
		if (write_en==1'b1)
			r_53_13 <= data_in;
	if (addr_selector[53]&addr_selector[14])
		data_out <= r_53_14;
		if (write_en==1'b1)
			r_53_14 <= data_in;
	if (addr_selector[53]&addr_selector[15])
		data_out <= r_53_15;
		if (write_en==1'b1)
			r_53_15 <= data_in;
	if (addr_selector[53]&addr_selector[16])
		data_out <= r_53_16;
		if (write_en==1'b1)
			r_53_16 <= data_in;
	if (addr_selector[53]&addr_selector[17])
		data_out <= r_53_17;
		if (write_en==1'b1)
			r_53_17 <= data_in;
	if (addr_selector[53]&addr_selector[18])
		data_out <= r_53_18;
		if (write_en==1'b1)
			r_53_18 <= data_in;
	if (addr_selector[53]&addr_selector[19])
		data_out <= r_53_19;
		if (write_en==1'b1)
			r_53_19 <= data_in;
	if (addr_selector[53]&addr_selector[20])
		data_out <= r_53_20;
		if (write_en==1'b1)
			r_53_20 <= data_in;
	if (addr_selector[53]&addr_selector[21])
		data_out <= r_53_21;
		if (write_en==1'b1)
			r_53_21 <= data_in;
	if (addr_selector[53]&addr_selector[22])
		data_out <= r_53_22;
		if (write_en==1'b1)
			r_53_22 <= data_in;
	if (addr_selector[53]&addr_selector[23])
		data_out <= r_53_23;
		if (write_en==1'b1)
			r_53_23 <= data_in;
	if (addr_selector[53]&addr_selector[24])
		data_out <= r_53_24;
		if (write_en==1'b1)
			r_53_24 <= data_in;
	if (addr_selector[53]&addr_selector[25])
		data_out <= r_53_25;
		if (write_en==1'b1)
			r_53_25 <= data_in;
	if (addr_selector[53]&addr_selector[26])
		data_out <= r_53_26;
		if (write_en==1'b1)
			r_53_26 <= data_in;
	if (addr_selector[53]&addr_selector[27])
		data_out <= r_53_27;
		if (write_en==1'b1)
			r_53_27 <= data_in;
	if (addr_selector[53]&addr_selector[28])
		data_out <= r_53_28;
		if (write_en==1'b1)
			r_53_28 <= data_in;
	if (addr_selector[53]&addr_selector[29])
		data_out <= r_53_29;
		if (write_en==1'b1)
			r_53_29 <= data_in;
	if (addr_selector[53]&addr_selector[30])
		data_out <= r_53_30;
		if (write_en==1'b1)
			r_53_30 <= data_in;
	if (addr_selector[53]&addr_selector[31])
		data_out <= r_53_31;
		if (write_en==1'b1)
			r_53_31 <= data_in;
	if (addr_selector[53]&addr_selector[32])
		data_out <= r_53_32;
		if (write_en==1'b1)
			r_53_32 <= data_in;
	if (addr_selector[53]&addr_selector[33])
		data_out <= r_53_33;
		if (write_en==1'b1)
			r_53_33 <= data_in;
	if (addr_selector[53]&addr_selector[34])
		data_out <= r_53_34;
		if (write_en==1'b1)
			r_53_34 <= data_in;
	if (addr_selector[53]&addr_selector[35])
		data_out <= r_53_35;
		if (write_en==1'b1)
			r_53_35 <= data_in;
	if (addr_selector[53]&addr_selector[36])
		data_out <= r_53_36;
		if (write_en==1'b1)
			r_53_36 <= data_in;
	if (addr_selector[53]&addr_selector[37])
		data_out <= r_53_37;
		if (write_en==1'b1)
			r_53_37 <= data_in;
	if (addr_selector[53]&addr_selector[38])
		data_out <= r_53_38;
		if (write_en==1'b1)
			r_53_38 <= data_in;
	if (addr_selector[53]&addr_selector[39])
		data_out <= r_53_39;
		if (write_en==1'b1)
			r_53_39 <= data_in;
	if (addr_selector[53]&addr_selector[40])
		data_out <= r_53_40;
		if (write_en==1'b1)
			r_53_40 <= data_in;
	if (addr_selector[53]&addr_selector[41])
		data_out <= r_53_41;
		if (write_en==1'b1)
			r_53_41 <= data_in;
	if (addr_selector[53]&addr_selector[42])
		data_out <= r_53_42;
		if (write_en==1'b1)
			r_53_42 <= data_in;
	if (addr_selector[53]&addr_selector[43])
		data_out <= r_53_43;
		if (write_en==1'b1)
			r_53_43 <= data_in;
	if (addr_selector[53]&addr_selector[44])
		data_out <= r_53_44;
		if (write_en==1'b1)
			r_53_44 <= data_in;
	if (addr_selector[53]&addr_selector[45])
		data_out <= r_53_45;
		if (write_en==1'b1)
			r_53_45 <= data_in;
	if (addr_selector[53]&addr_selector[46])
		data_out <= r_53_46;
		if (write_en==1'b1)
			r_53_46 <= data_in;
	if (addr_selector[53]&addr_selector[47])
		data_out <= r_53_47;
		if (write_en==1'b1)
			r_53_47 <= data_in;
	if (addr_selector[53]&addr_selector[48])
		data_out <= r_53_48;
		if (write_en==1'b1)
			r_53_48 <= data_in;
	if (addr_selector[53]&addr_selector[49])
		data_out <= r_53_49;
		if (write_en==1'b1)
			r_53_49 <= data_in;
	if (addr_selector[53]&addr_selector[50])
		data_out <= r_53_50;
		if (write_en==1'b1)
			r_53_50 <= data_in;
	if (addr_selector[53]&addr_selector[51])
		data_out <= r_53_51;
		if (write_en==1'b1)
			r_53_51 <= data_in;
	if (addr_selector[53]&addr_selector[52])
		data_out <= r_53_52;
		if (write_en==1'b1)
			r_53_52 <= data_in;
	if (addr_selector[53]&addr_selector[53])
		data_out <= r_53_53;
		if (write_en==1'b1)
			r_53_53 <= data_in;
	if (addr_selector[53]&addr_selector[54])
		data_out <= r_53_54;
		if (write_en==1'b1)
			r_53_54 <= data_in;
	if (addr_selector[53]&addr_selector[55])
		data_out <= r_53_55;
		if (write_en==1'b1)
			r_53_55 <= data_in;
	if (addr_selector[53]&addr_selector[56])
		data_out <= r_53_56;
		if (write_en==1'b1)
			r_53_56 <= data_in;
	if (addr_selector[53]&addr_selector[57])
		data_out <= r_53_57;
		if (write_en==1'b1)
			r_53_57 <= data_in;
	if (addr_selector[53]&addr_selector[58])
		data_out <= r_53_58;
		if (write_en==1'b1)
			r_53_58 <= data_in;
	if (addr_selector[53]&addr_selector[59])
		data_out <= r_53_59;
		if (write_en==1'b1)
			r_53_59 <= data_in;
	if (addr_selector[53]&addr_selector[60])
		data_out <= r_53_60;
		if (write_en==1'b1)
			r_53_60 <= data_in;
	if (addr_selector[53]&addr_selector[61])
		data_out <= r_53_61;
		if (write_en==1'b1)
			r_53_61 <= data_in;
	if (addr_selector[53]&addr_selector[62])
		data_out <= r_53_62;
		if (write_en==1'b1)
			r_53_62 <= data_in;
	if (addr_selector[53]&addr_selector[63])
		data_out <= r_53_63;
		if (write_en==1'b1)
			r_53_63 <= data_in;
	if (addr_selector[54]&addr_selector[0])
		data_out <= r_54_0;
		if (write_en==1'b1)
			r_54_0 <= data_in;
	if (addr_selector[54]&addr_selector[1])
		data_out <= r_54_1;
		if (write_en==1'b1)
			r_54_1 <= data_in;
	if (addr_selector[54]&addr_selector[2])
		data_out <= r_54_2;
		if (write_en==1'b1)
			r_54_2 <= data_in;
	if (addr_selector[54]&addr_selector[3])
		data_out <= r_54_3;
		if (write_en==1'b1)
			r_54_3 <= data_in;
	if (addr_selector[54]&addr_selector[4])
		data_out <= r_54_4;
		if (write_en==1'b1)
			r_54_4 <= data_in;
	if (addr_selector[54]&addr_selector[5])
		data_out <= r_54_5;
		if (write_en==1'b1)
			r_54_5 <= data_in;
	if (addr_selector[54]&addr_selector[6])
		data_out <= r_54_6;
		if (write_en==1'b1)
			r_54_6 <= data_in;
	if (addr_selector[54]&addr_selector[7])
		data_out <= r_54_7;
		if (write_en==1'b1)
			r_54_7 <= data_in;
	if (addr_selector[54]&addr_selector[8])
		data_out <= r_54_8;
		if (write_en==1'b1)
			r_54_8 <= data_in;
	if (addr_selector[54]&addr_selector[9])
		data_out <= r_54_9;
		if (write_en==1'b1)
			r_54_9 <= data_in;
	if (addr_selector[54]&addr_selector[10])
		data_out <= r_54_10;
		if (write_en==1'b1)
			r_54_10 <= data_in;
	if (addr_selector[54]&addr_selector[11])
		data_out <= r_54_11;
		if (write_en==1'b1)
			r_54_11 <= data_in;
	if (addr_selector[54]&addr_selector[12])
		data_out <= r_54_12;
		if (write_en==1'b1)
			r_54_12 <= data_in;
	if (addr_selector[54]&addr_selector[13])
		data_out <= r_54_13;
		if (write_en==1'b1)
			r_54_13 <= data_in;
	if (addr_selector[54]&addr_selector[14])
		data_out <= r_54_14;
		if (write_en==1'b1)
			r_54_14 <= data_in;
	if (addr_selector[54]&addr_selector[15])
		data_out <= r_54_15;
		if (write_en==1'b1)
			r_54_15 <= data_in;
	if (addr_selector[54]&addr_selector[16])
		data_out <= r_54_16;
		if (write_en==1'b1)
			r_54_16 <= data_in;
	if (addr_selector[54]&addr_selector[17])
		data_out <= r_54_17;
		if (write_en==1'b1)
			r_54_17 <= data_in;
	if (addr_selector[54]&addr_selector[18])
		data_out <= r_54_18;
		if (write_en==1'b1)
			r_54_18 <= data_in;
	if (addr_selector[54]&addr_selector[19])
		data_out <= r_54_19;
		if (write_en==1'b1)
			r_54_19 <= data_in;
	if (addr_selector[54]&addr_selector[20])
		data_out <= r_54_20;
		if (write_en==1'b1)
			r_54_20 <= data_in;
	if (addr_selector[54]&addr_selector[21])
		data_out <= r_54_21;
		if (write_en==1'b1)
			r_54_21 <= data_in;
	if (addr_selector[54]&addr_selector[22])
		data_out <= r_54_22;
		if (write_en==1'b1)
			r_54_22 <= data_in;
	if (addr_selector[54]&addr_selector[23])
		data_out <= r_54_23;
		if (write_en==1'b1)
			r_54_23 <= data_in;
	if (addr_selector[54]&addr_selector[24])
		data_out <= r_54_24;
		if (write_en==1'b1)
			r_54_24 <= data_in;
	if (addr_selector[54]&addr_selector[25])
		data_out <= r_54_25;
		if (write_en==1'b1)
			r_54_25 <= data_in;
	if (addr_selector[54]&addr_selector[26])
		data_out <= r_54_26;
		if (write_en==1'b1)
			r_54_26 <= data_in;
	if (addr_selector[54]&addr_selector[27])
		data_out <= r_54_27;
		if (write_en==1'b1)
			r_54_27 <= data_in;
	if (addr_selector[54]&addr_selector[28])
		data_out <= r_54_28;
		if (write_en==1'b1)
			r_54_28 <= data_in;
	if (addr_selector[54]&addr_selector[29])
		data_out <= r_54_29;
		if (write_en==1'b1)
			r_54_29 <= data_in;
	if (addr_selector[54]&addr_selector[30])
		data_out <= r_54_30;
		if (write_en==1'b1)
			r_54_30 <= data_in;
	if (addr_selector[54]&addr_selector[31])
		data_out <= r_54_31;
		if (write_en==1'b1)
			r_54_31 <= data_in;
	if (addr_selector[54]&addr_selector[32])
		data_out <= r_54_32;
		if (write_en==1'b1)
			r_54_32 <= data_in;
	if (addr_selector[54]&addr_selector[33])
		data_out <= r_54_33;
		if (write_en==1'b1)
			r_54_33 <= data_in;
	if (addr_selector[54]&addr_selector[34])
		data_out <= r_54_34;
		if (write_en==1'b1)
			r_54_34 <= data_in;
	if (addr_selector[54]&addr_selector[35])
		data_out <= r_54_35;
		if (write_en==1'b1)
			r_54_35 <= data_in;
	if (addr_selector[54]&addr_selector[36])
		data_out <= r_54_36;
		if (write_en==1'b1)
			r_54_36 <= data_in;
	if (addr_selector[54]&addr_selector[37])
		data_out <= r_54_37;
		if (write_en==1'b1)
			r_54_37 <= data_in;
	if (addr_selector[54]&addr_selector[38])
		data_out <= r_54_38;
		if (write_en==1'b1)
			r_54_38 <= data_in;
	if (addr_selector[54]&addr_selector[39])
		data_out <= r_54_39;
		if (write_en==1'b1)
			r_54_39 <= data_in;
	if (addr_selector[54]&addr_selector[40])
		data_out <= r_54_40;
		if (write_en==1'b1)
			r_54_40 <= data_in;
	if (addr_selector[54]&addr_selector[41])
		data_out <= r_54_41;
		if (write_en==1'b1)
			r_54_41 <= data_in;
	if (addr_selector[54]&addr_selector[42])
		data_out <= r_54_42;
		if (write_en==1'b1)
			r_54_42 <= data_in;
	if (addr_selector[54]&addr_selector[43])
		data_out <= r_54_43;
		if (write_en==1'b1)
			r_54_43 <= data_in;
	if (addr_selector[54]&addr_selector[44])
		data_out <= r_54_44;
		if (write_en==1'b1)
			r_54_44 <= data_in;
	if (addr_selector[54]&addr_selector[45])
		data_out <= r_54_45;
		if (write_en==1'b1)
			r_54_45 <= data_in;
	if (addr_selector[54]&addr_selector[46])
		data_out <= r_54_46;
		if (write_en==1'b1)
			r_54_46 <= data_in;
	if (addr_selector[54]&addr_selector[47])
		data_out <= r_54_47;
		if (write_en==1'b1)
			r_54_47 <= data_in;
	if (addr_selector[54]&addr_selector[48])
		data_out <= r_54_48;
		if (write_en==1'b1)
			r_54_48 <= data_in;
	if (addr_selector[54]&addr_selector[49])
		data_out <= r_54_49;
		if (write_en==1'b1)
			r_54_49 <= data_in;
	if (addr_selector[54]&addr_selector[50])
		data_out <= r_54_50;
		if (write_en==1'b1)
			r_54_50 <= data_in;
	if (addr_selector[54]&addr_selector[51])
		data_out <= r_54_51;
		if (write_en==1'b1)
			r_54_51 <= data_in;
	if (addr_selector[54]&addr_selector[52])
		data_out <= r_54_52;
		if (write_en==1'b1)
			r_54_52 <= data_in;
	if (addr_selector[54]&addr_selector[53])
		data_out <= r_54_53;
		if (write_en==1'b1)
			r_54_53 <= data_in;
	if (addr_selector[54]&addr_selector[54])
		data_out <= r_54_54;
		if (write_en==1'b1)
			r_54_54 <= data_in;
	if (addr_selector[54]&addr_selector[55])
		data_out <= r_54_55;
		if (write_en==1'b1)
			r_54_55 <= data_in;
	if (addr_selector[54]&addr_selector[56])
		data_out <= r_54_56;
		if (write_en==1'b1)
			r_54_56 <= data_in;
	if (addr_selector[54]&addr_selector[57])
		data_out <= r_54_57;
		if (write_en==1'b1)
			r_54_57 <= data_in;
	if (addr_selector[54]&addr_selector[58])
		data_out <= r_54_58;
		if (write_en==1'b1)
			r_54_58 <= data_in;
	if (addr_selector[54]&addr_selector[59])
		data_out <= r_54_59;
		if (write_en==1'b1)
			r_54_59 <= data_in;
	if (addr_selector[54]&addr_selector[60])
		data_out <= r_54_60;
		if (write_en==1'b1)
			r_54_60 <= data_in;
	if (addr_selector[54]&addr_selector[61])
		data_out <= r_54_61;
		if (write_en==1'b1)
			r_54_61 <= data_in;
	if (addr_selector[54]&addr_selector[62])
		data_out <= r_54_62;
		if (write_en==1'b1)
			r_54_62 <= data_in;
	if (addr_selector[54]&addr_selector[63])
		data_out <= r_54_63;
		if (write_en==1'b1)
			r_54_63 <= data_in;
	if (addr_selector[55]&addr_selector[0])
		data_out <= r_55_0;
		if (write_en==1'b1)
			r_55_0 <= data_in;
	if (addr_selector[55]&addr_selector[1])
		data_out <= r_55_1;
		if (write_en==1'b1)
			r_55_1 <= data_in;
	if (addr_selector[55]&addr_selector[2])
		data_out <= r_55_2;
		if (write_en==1'b1)
			r_55_2 <= data_in;
	if (addr_selector[55]&addr_selector[3])
		data_out <= r_55_3;
		if (write_en==1'b1)
			r_55_3 <= data_in;
	if (addr_selector[55]&addr_selector[4])
		data_out <= r_55_4;
		if (write_en==1'b1)
			r_55_4 <= data_in;
	if (addr_selector[55]&addr_selector[5])
		data_out <= r_55_5;
		if (write_en==1'b1)
			r_55_5 <= data_in;
	if (addr_selector[55]&addr_selector[6])
		data_out <= r_55_6;
		if (write_en==1'b1)
			r_55_6 <= data_in;
	if (addr_selector[55]&addr_selector[7])
		data_out <= r_55_7;
		if (write_en==1'b1)
			r_55_7 <= data_in;
	if (addr_selector[55]&addr_selector[8])
		data_out <= r_55_8;
		if (write_en==1'b1)
			r_55_8 <= data_in;
	if (addr_selector[55]&addr_selector[9])
		data_out <= r_55_9;
		if (write_en==1'b1)
			r_55_9 <= data_in;
	if (addr_selector[55]&addr_selector[10])
		data_out <= r_55_10;
		if (write_en==1'b1)
			r_55_10 <= data_in;
	if (addr_selector[55]&addr_selector[11])
		data_out <= r_55_11;
		if (write_en==1'b1)
			r_55_11 <= data_in;
	if (addr_selector[55]&addr_selector[12])
		data_out <= r_55_12;
		if (write_en==1'b1)
			r_55_12 <= data_in;
	if (addr_selector[55]&addr_selector[13])
		data_out <= r_55_13;
		if (write_en==1'b1)
			r_55_13 <= data_in;
	if (addr_selector[55]&addr_selector[14])
		data_out <= r_55_14;
		if (write_en==1'b1)
			r_55_14 <= data_in;
	if (addr_selector[55]&addr_selector[15])
		data_out <= r_55_15;
		if (write_en==1'b1)
			r_55_15 <= data_in;
	if (addr_selector[55]&addr_selector[16])
		data_out <= r_55_16;
		if (write_en==1'b1)
			r_55_16 <= data_in;
	if (addr_selector[55]&addr_selector[17])
		data_out <= r_55_17;
		if (write_en==1'b1)
			r_55_17 <= data_in;
	if (addr_selector[55]&addr_selector[18])
		data_out <= r_55_18;
		if (write_en==1'b1)
			r_55_18 <= data_in;
	if (addr_selector[55]&addr_selector[19])
		data_out <= r_55_19;
		if (write_en==1'b1)
			r_55_19 <= data_in;
	if (addr_selector[55]&addr_selector[20])
		data_out <= r_55_20;
		if (write_en==1'b1)
			r_55_20 <= data_in;
	if (addr_selector[55]&addr_selector[21])
		data_out <= r_55_21;
		if (write_en==1'b1)
			r_55_21 <= data_in;
	if (addr_selector[55]&addr_selector[22])
		data_out <= r_55_22;
		if (write_en==1'b1)
			r_55_22 <= data_in;
	if (addr_selector[55]&addr_selector[23])
		data_out <= r_55_23;
		if (write_en==1'b1)
			r_55_23 <= data_in;
	if (addr_selector[55]&addr_selector[24])
		data_out <= r_55_24;
		if (write_en==1'b1)
			r_55_24 <= data_in;
	if (addr_selector[55]&addr_selector[25])
		data_out <= r_55_25;
		if (write_en==1'b1)
			r_55_25 <= data_in;
	if (addr_selector[55]&addr_selector[26])
		data_out <= r_55_26;
		if (write_en==1'b1)
			r_55_26 <= data_in;
	if (addr_selector[55]&addr_selector[27])
		data_out <= r_55_27;
		if (write_en==1'b1)
			r_55_27 <= data_in;
	if (addr_selector[55]&addr_selector[28])
		data_out <= r_55_28;
		if (write_en==1'b1)
			r_55_28 <= data_in;
	if (addr_selector[55]&addr_selector[29])
		data_out <= r_55_29;
		if (write_en==1'b1)
			r_55_29 <= data_in;
	if (addr_selector[55]&addr_selector[30])
		data_out <= r_55_30;
		if (write_en==1'b1)
			r_55_30 <= data_in;
	if (addr_selector[55]&addr_selector[31])
		data_out <= r_55_31;
		if (write_en==1'b1)
			r_55_31 <= data_in;
	if (addr_selector[55]&addr_selector[32])
		data_out <= r_55_32;
		if (write_en==1'b1)
			r_55_32 <= data_in;
	if (addr_selector[55]&addr_selector[33])
		data_out <= r_55_33;
		if (write_en==1'b1)
			r_55_33 <= data_in;
	if (addr_selector[55]&addr_selector[34])
		data_out <= r_55_34;
		if (write_en==1'b1)
			r_55_34 <= data_in;
	if (addr_selector[55]&addr_selector[35])
		data_out <= r_55_35;
		if (write_en==1'b1)
			r_55_35 <= data_in;
	if (addr_selector[55]&addr_selector[36])
		data_out <= r_55_36;
		if (write_en==1'b1)
			r_55_36 <= data_in;
	if (addr_selector[55]&addr_selector[37])
		data_out <= r_55_37;
		if (write_en==1'b1)
			r_55_37 <= data_in;
	if (addr_selector[55]&addr_selector[38])
		data_out <= r_55_38;
		if (write_en==1'b1)
			r_55_38 <= data_in;
	if (addr_selector[55]&addr_selector[39])
		data_out <= r_55_39;
		if (write_en==1'b1)
			r_55_39 <= data_in;
	if (addr_selector[55]&addr_selector[40])
		data_out <= r_55_40;
		if (write_en==1'b1)
			r_55_40 <= data_in;
	if (addr_selector[55]&addr_selector[41])
		data_out <= r_55_41;
		if (write_en==1'b1)
			r_55_41 <= data_in;
	if (addr_selector[55]&addr_selector[42])
		data_out <= r_55_42;
		if (write_en==1'b1)
			r_55_42 <= data_in;
	if (addr_selector[55]&addr_selector[43])
		data_out <= r_55_43;
		if (write_en==1'b1)
			r_55_43 <= data_in;
	if (addr_selector[55]&addr_selector[44])
		data_out <= r_55_44;
		if (write_en==1'b1)
			r_55_44 <= data_in;
	if (addr_selector[55]&addr_selector[45])
		data_out <= r_55_45;
		if (write_en==1'b1)
			r_55_45 <= data_in;
	if (addr_selector[55]&addr_selector[46])
		data_out <= r_55_46;
		if (write_en==1'b1)
			r_55_46 <= data_in;
	if (addr_selector[55]&addr_selector[47])
		data_out <= r_55_47;
		if (write_en==1'b1)
			r_55_47 <= data_in;
	if (addr_selector[55]&addr_selector[48])
		data_out <= r_55_48;
		if (write_en==1'b1)
			r_55_48 <= data_in;
	if (addr_selector[55]&addr_selector[49])
		data_out <= r_55_49;
		if (write_en==1'b1)
			r_55_49 <= data_in;
	if (addr_selector[55]&addr_selector[50])
		data_out <= r_55_50;
		if (write_en==1'b1)
			r_55_50 <= data_in;
	if (addr_selector[55]&addr_selector[51])
		data_out <= r_55_51;
		if (write_en==1'b1)
			r_55_51 <= data_in;
	if (addr_selector[55]&addr_selector[52])
		data_out <= r_55_52;
		if (write_en==1'b1)
			r_55_52 <= data_in;
	if (addr_selector[55]&addr_selector[53])
		data_out <= r_55_53;
		if (write_en==1'b1)
			r_55_53 <= data_in;
	if (addr_selector[55]&addr_selector[54])
		data_out <= r_55_54;
		if (write_en==1'b1)
			r_55_54 <= data_in;
	if (addr_selector[55]&addr_selector[55])
		data_out <= r_55_55;
		if (write_en==1'b1)
			r_55_55 <= data_in;
	if (addr_selector[55]&addr_selector[56])
		data_out <= r_55_56;
		if (write_en==1'b1)
			r_55_56 <= data_in;
	if (addr_selector[55]&addr_selector[57])
		data_out <= r_55_57;
		if (write_en==1'b1)
			r_55_57 <= data_in;
	if (addr_selector[55]&addr_selector[58])
		data_out <= r_55_58;
		if (write_en==1'b1)
			r_55_58 <= data_in;
	if (addr_selector[55]&addr_selector[59])
		data_out <= r_55_59;
		if (write_en==1'b1)
			r_55_59 <= data_in;
	if (addr_selector[55]&addr_selector[60])
		data_out <= r_55_60;
		if (write_en==1'b1)
			r_55_60 <= data_in;
	if (addr_selector[55]&addr_selector[61])
		data_out <= r_55_61;
		if (write_en==1'b1)
			r_55_61 <= data_in;
	if (addr_selector[55]&addr_selector[62])
		data_out <= r_55_62;
		if (write_en==1'b1)
			r_55_62 <= data_in;
	if (addr_selector[55]&addr_selector[63])
		data_out <= r_55_63;
		if (write_en==1'b1)
			r_55_63 <= data_in;
	if (addr_selector[56]&addr_selector[0])
		data_out <= r_56_0;
		if (write_en==1'b1)
			r_56_0 <= data_in;
	if (addr_selector[56]&addr_selector[1])
		data_out <= r_56_1;
		if (write_en==1'b1)
			r_56_1 <= data_in;
	if (addr_selector[56]&addr_selector[2])
		data_out <= r_56_2;
		if (write_en==1'b1)
			r_56_2 <= data_in;
	if (addr_selector[56]&addr_selector[3])
		data_out <= r_56_3;
		if (write_en==1'b1)
			r_56_3 <= data_in;
	if (addr_selector[56]&addr_selector[4])
		data_out <= r_56_4;
		if (write_en==1'b1)
			r_56_4 <= data_in;
	if (addr_selector[56]&addr_selector[5])
		data_out <= r_56_5;
		if (write_en==1'b1)
			r_56_5 <= data_in;
	if (addr_selector[56]&addr_selector[6])
		data_out <= r_56_6;
		if (write_en==1'b1)
			r_56_6 <= data_in;
	if (addr_selector[56]&addr_selector[7])
		data_out <= r_56_7;
		if (write_en==1'b1)
			r_56_7 <= data_in;
	if (addr_selector[56]&addr_selector[8])
		data_out <= r_56_8;
		if (write_en==1'b1)
			r_56_8 <= data_in;
	if (addr_selector[56]&addr_selector[9])
		data_out <= r_56_9;
		if (write_en==1'b1)
			r_56_9 <= data_in;
	if (addr_selector[56]&addr_selector[10])
		data_out <= r_56_10;
		if (write_en==1'b1)
			r_56_10 <= data_in;
	if (addr_selector[56]&addr_selector[11])
		data_out <= r_56_11;
		if (write_en==1'b1)
			r_56_11 <= data_in;
	if (addr_selector[56]&addr_selector[12])
		data_out <= r_56_12;
		if (write_en==1'b1)
			r_56_12 <= data_in;
	if (addr_selector[56]&addr_selector[13])
		data_out <= r_56_13;
		if (write_en==1'b1)
			r_56_13 <= data_in;
	if (addr_selector[56]&addr_selector[14])
		data_out <= r_56_14;
		if (write_en==1'b1)
			r_56_14 <= data_in;
	if (addr_selector[56]&addr_selector[15])
		data_out <= r_56_15;
		if (write_en==1'b1)
			r_56_15 <= data_in;
	if (addr_selector[56]&addr_selector[16])
		data_out <= r_56_16;
		if (write_en==1'b1)
			r_56_16 <= data_in;
	if (addr_selector[56]&addr_selector[17])
		data_out <= r_56_17;
		if (write_en==1'b1)
			r_56_17 <= data_in;
	if (addr_selector[56]&addr_selector[18])
		data_out <= r_56_18;
		if (write_en==1'b1)
			r_56_18 <= data_in;
	if (addr_selector[56]&addr_selector[19])
		data_out <= r_56_19;
		if (write_en==1'b1)
			r_56_19 <= data_in;
	if (addr_selector[56]&addr_selector[20])
		data_out <= r_56_20;
		if (write_en==1'b1)
			r_56_20 <= data_in;
	if (addr_selector[56]&addr_selector[21])
		data_out <= r_56_21;
		if (write_en==1'b1)
			r_56_21 <= data_in;
	if (addr_selector[56]&addr_selector[22])
		data_out <= r_56_22;
		if (write_en==1'b1)
			r_56_22 <= data_in;
	if (addr_selector[56]&addr_selector[23])
		data_out <= r_56_23;
		if (write_en==1'b1)
			r_56_23 <= data_in;
	if (addr_selector[56]&addr_selector[24])
		data_out <= r_56_24;
		if (write_en==1'b1)
			r_56_24 <= data_in;
	if (addr_selector[56]&addr_selector[25])
		data_out <= r_56_25;
		if (write_en==1'b1)
			r_56_25 <= data_in;
	if (addr_selector[56]&addr_selector[26])
		data_out <= r_56_26;
		if (write_en==1'b1)
			r_56_26 <= data_in;
	if (addr_selector[56]&addr_selector[27])
		data_out <= r_56_27;
		if (write_en==1'b1)
			r_56_27 <= data_in;
	if (addr_selector[56]&addr_selector[28])
		data_out <= r_56_28;
		if (write_en==1'b1)
			r_56_28 <= data_in;
	if (addr_selector[56]&addr_selector[29])
		data_out <= r_56_29;
		if (write_en==1'b1)
			r_56_29 <= data_in;
	if (addr_selector[56]&addr_selector[30])
		data_out <= r_56_30;
		if (write_en==1'b1)
			r_56_30 <= data_in;
	if (addr_selector[56]&addr_selector[31])
		data_out <= r_56_31;
		if (write_en==1'b1)
			r_56_31 <= data_in;
	if (addr_selector[56]&addr_selector[32])
		data_out <= r_56_32;
		if (write_en==1'b1)
			r_56_32 <= data_in;
	if (addr_selector[56]&addr_selector[33])
		data_out <= r_56_33;
		if (write_en==1'b1)
			r_56_33 <= data_in;
	if (addr_selector[56]&addr_selector[34])
		data_out <= r_56_34;
		if (write_en==1'b1)
			r_56_34 <= data_in;
	if (addr_selector[56]&addr_selector[35])
		data_out <= r_56_35;
		if (write_en==1'b1)
			r_56_35 <= data_in;
	if (addr_selector[56]&addr_selector[36])
		data_out <= r_56_36;
		if (write_en==1'b1)
			r_56_36 <= data_in;
	if (addr_selector[56]&addr_selector[37])
		data_out <= r_56_37;
		if (write_en==1'b1)
			r_56_37 <= data_in;
	if (addr_selector[56]&addr_selector[38])
		data_out <= r_56_38;
		if (write_en==1'b1)
			r_56_38 <= data_in;
	if (addr_selector[56]&addr_selector[39])
		data_out <= r_56_39;
		if (write_en==1'b1)
			r_56_39 <= data_in;
	if (addr_selector[56]&addr_selector[40])
		data_out <= r_56_40;
		if (write_en==1'b1)
			r_56_40 <= data_in;
	if (addr_selector[56]&addr_selector[41])
		data_out <= r_56_41;
		if (write_en==1'b1)
			r_56_41 <= data_in;
	if (addr_selector[56]&addr_selector[42])
		data_out <= r_56_42;
		if (write_en==1'b1)
			r_56_42 <= data_in;
	if (addr_selector[56]&addr_selector[43])
		data_out <= r_56_43;
		if (write_en==1'b1)
			r_56_43 <= data_in;
	if (addr_selector[56]&addr_selector[44])
		data_out <= r_56_44;
		if (write_en==1'b1)
			r_56_44 <= data_in;
	if (addr_selector[56]&addr_selector[45])
		data_out <= r_56_45;
		if (write_en==1'b1)
			r_56_45 <= data_in;
	if (addr_selector[56]&addr_selector[46])
		data_out <= r_56_46;
		if (write_en==1'b1)
			r_56_46 <= data_in;
	if (addr_selector[56]&addr_selector[47])
		data_out <= r_56_47;
		if (write_en==1'b1)
			r_56_47 <= data_in;
	if (addr_selector[56]&addr_selector[48])
		data_out <= r_56_48;
		if (write_en==1'b1)
			r_56_48 <= data_in;
	if (addr_selector[56]&addr_selector[49])
		data_out <= r_56_49;
		if (write_en==1'b1)
			r_56_49 <= data_in;
	if (addr_selector[56]&addr_selector[50])
		data_out <= r_56_50;
		if (write_en==1'b1)
			r_56_50 <= data_in;
	if (addr_selector[56]&addr_selector[51])
		data_out <= r_56_51;
		if (write_en==1'b1)
			r_56_51 <= data_in;
	if (addr_selector[56]&addr_selector[52])
		data_out <= r_56_52;
		if (write_en==1'b1)
			r_56_52 <= data_in;
	if (addr_selector[56]&addr_selector[53])
		data_out <= r_56_53;
		if (write_en==1'b1)
			r_56_53 <= data_in;
	if (addr_selector[56]&addr_selector[54])
		data_out <= r_56_54;
		if (write_en==1'b1)
			r_56_54 <= data_in;
	if (addr_selector[56]&addr_selector[55])
		data_out <= r_56_55;
		if (write_en==1'b1)
			r_56_55 <= data_in;
	if (addr_selector[56]&addr_selector[56])
		data_out <= r_56_56;
		if (write_en==1'b1)
			r_56_56 <= data_in;
	if (addr_selector[56]&addr_selector[57])
		data_out <= r_56_57;
		if (write_en==1'b1)
			r_56_57 <= data_in;
	if (addr_selector[56]&addr_selector[58])
		data_out <= r_56_58;
		if (write_en==1'b1)
			r_56_58 <= data_in;
	if (addr_selector[56]&addr_selector[59])
		data_out <= r_56_59;
		if (write_en==1'b1)
			r_56_59 <= data_in;
	if (addr_selector[56]&addr_selector[60])
		data_out <= r_56_60;
		if (write_en==1'b1)
			r_56_60 <= data_in;
	if (addr_selector[56]&addr_selector[61])
		data_out <= r_56_61;
		if (write_en==1'b1)
			r_56_61 <= data_in;
	if (addr_selector[56]&addr_selector[62])
		data_out <= r_56_62;
		if (write_en==1'b1)
			r_56_62 <= data_in;
	if (addr_selector[56]&addr_selector[63])
		data_out <= r_56_63;
		if (write_en==1'b1)
			r_56_63 <= data_in;
	if (addr_selector[57]&addr_selector[0])
		data_out <= r_57_0;
		if (write_en==1'b1)
			r_57_0 <= data_in;
	if (addr_selector[57]&addr_selector[1])
		data_out <= r_57_1;
		if (write_en==1'b1)
			r_57_1 <= data_in;
	if (addr_selector[57]&addr_selector[2])
		data_out <= r_57_2;
		if (write_en==1'b1)
			r_57_2 <= data_in;
	if (addr_selector[57]&addr_selector[3])
		data_out <= r_57_3;
		if (write_en==1'b1)
			r_57_3 <= data_in;
	if (addr_selector[57]&addr_selector[4])
		data_out <= r_57_4;
		if (write_en==1'b1)
			r_57_4 <= data_in;
	if (addr_selector[57]&addr_selector[5])
		data_out <= r_57_5;
		if (write_en==1'b1)
			r_57_5 <= data_in;
	if (addr_selector[57]&addr_selector[6])
		data_out <= r_57_6;
		if (write_en==1'b1)
			r_57_6 <= data_in;
	if (addr_selector[57]&addr_selector[7])
		data_out <= r_57_7;
		if (write_en==1'b1)
			r_57_7 <= data_in;
	if (addr_selector[57]&addr_selector[8])
		data_out <= r_57_8;
		if (write_en==1'b1)
			r_57_8 <= data_in;
	if (addr_selector[57]&addr_selector[9])
		data_out <= r_57_9;
		if (write_en==1'b1)
			r_57_9 <= data_in;
	if (addr_selector[57]&addr_selector[10])
		data_out <= r_57_10;
		if (write_en==1'b1)
			r_57_10 <= data_in;
	if (addr_selector[57]&addr_selector[11])
		data_out <= r_57_11;
		if (write_en==1'b1)
			r_57_11 <= data_in;
	if (addr_selector[57]&addr_selector[12])
		data_out <= r_57_12;
		if (write_en==1'b1)
			r_57_12 <= data_in;
	if (addr_selector[57]&addr_selector[13])
		data_out <= r_57_13;
		if (write_en==1'b1)
			r_57_13 <= data_in;
	if (addr_selector[57]&addr_selector[14])
		data_out <= r_57_14;
		if (write_en==1'b1)
			r_57_14 <= data_in;
	if (addr_selector[57]&addr_selector[15])
		data_out <= r_57_15;
		if (write_en==1'b1)
			r_57_15 <= data_in;
	if (addr_selector[57]&addr_selector[16])
		data_out <= r_57_16;
		if (write_en==1'b1)
			r_57_16 <= data_in;
	if (addr_selector[57]&addr_selector[17])
		data_out <= r_57_17;
		if (write_en==1'b1)
			r_57_17 <= data_in;
	if (addr_selector[57]&addr_selector[18])
		data_out <= r_57_18;
		if (write_en==1'b1)
			r_57_18 <= data_in;
	if (addr_selector[57]&addr_selector[19])
		data_out <= r_57_19;
		if (write_en==1'b1)
			r_57_19 <= data_in;
	if (addr_selector[57]&addr_selector[20])
		data_out <= r_57_20;
		if (write_en==1'b1)
			r_57_20 <= data_in;
	if (addr_selector[57]&addr_selector[21])
		data_out <= r_57_21;
		if (write_en==1'b1)
			r_57_21 <= data_in;
	if (addr_selector[57]&addr_selector[22])
		data_out <= r_57_22;
		if (write_en==1'b1)
			r_57_22 <= data_in;
	if (addr_selector[57]&addr_selector[23])
		data_out <= r_57_23;
		if (write_en==1'b1)
			r_57_23 <= data_in;
	if (addr_selector[57]&addr_selector[24])
		data_out <= r_57_24;
		if (write_en==1'b1)
			r_57_24 <= data_in;
	if (addr_selector[57]&addr_selector[25])
		data_out <= r_57_25;
		if (write_en==1'b1)
			r_57_25 <= data_in;
	if (addr_selector[57]&addr_selector[26])
		data_out <= r_57_26;
		if (write_en==1'b1)
			r_57_26 <= data_in;
	if (addr_selector[57]&addr_selector[27])
		data_out <= r_57_27;
		if (write_en==1'b1)
			r_57_27 <= data_in;
	if (addr_selector[57]&addr_selector[28])
		data_out <= r_57_28;
		if (write_en==1'b1)
			r_57_28 <= data_in;
	if (addr_selector[57]&addr_selector[29])
		data_out <= r_57_29;
		if (write_en==1'b1)
			r_57_29 <= data_in;
	if (addr_selector[57]&addr_selector[30])
		data_out <= r_57_30;
		if (write_en==1'b1)
			r_57_30 <= data_in;
	if (addr_selector[57]&addr_selector[31])
		data_out <= r_57_31;
		if (write_en==1'b1)
			r_57_31 <= data_in;
	if (addr_selector[57]&addr_selector[32])
		data_out <= r_57_32;
		if (write_en==1'b1)
			r_57_32 <= data_in;
	if (addr_selector[57]&addr_selector[33])
		data_out <= r_57_33;
		if (write_en==1'b1)
			r_57_33 <= data_in;
	if (addr_selector[57]&addr_selector[34])
		data_out <= r_57_34;
		if (write_en==1'b1)
			r_57_34 <= data_in;
	if (addr_selector[57]&addr_selector[35])
		data_out <= r_57_35;
		if (write_en==1'b1)
			r_57_35 <= data_in;
	if (addr_selector[57]&addr_selector[36])
		data_out <= r_57_36;
		if (write_en==1'b1)
			r_57_36 <= data_in;
	if (addr_selector[57]&addr_selector[37])
		data_out <= r_57_37;
		if (write_en==1'b1)
			r_57_37 <= data_in;
	if (addr_selector[57]&addr_selector[38])
		data_out <= r_57_38;
		if (write_en==1'b1)
			r_57_38 <= data_in;
	if (addr_selector[57]&addr_selector[39])
		data_out <= r_57_39;
		if (write_en==1'b1)
			r_57_39 <= data_in;
	if (addr_selector[57]&addr_selector[40])
		data_out <= r_57_40;
		if (write_en==1'b1)
			r_57_40 <= data_in;
	if (addr_selector[57]&addr_selector[41])
		data_out <= r_57_41;
		if (write_en==1'b1)
			r_57_41 <= data_in;
	if (addr_selector[57]&addr_selector[42])
		data_out <= r_57_42;
		if (write_en==1'b1)
			r_57_42 <= data_in;
	if (addr_selector[57]&addr_selector[43])
		data_out <= r_57_43;
		if (write_en==1'b1)
			r_57_43 <= data_in;
	if (addr_selector[57]&addr_selector[44])
		data_out <= r_57_44;
		if (write_en==1'b1)
			r_57_44 <= data_in;
	if (addr_selector[57]&addr_selector[45])
		data_out <= r_57_45;
		if (write_en==1'b1)
			r_57_45 <= data_in;
	if (addr_selector[57]&addr_selector[46])
		data_out <= r_57_46;
		if (write_en==1'b1)
			r_57_46 <= data_in;
	if (addr_selector[57]&addr_selector[47])
		data_out <= r_57_47;
		if (write_en==1'b1)
			r_57_47 <= data_in;
	if (addr_selector[57]&addr_selector[48])
		data_out <= r_57_48;
		if (write_en==1'b1)
			r_57_48 <= data_in;
	if (addr_selector[57]&addr_selector[49])
		data_out <= r_57_49;
		if (write_en==1'b1)
			r_57_49 <= data_in;
	if (addr_selector[57]&addr_selector[50])
		data_out <= r_57_50;
		if (write_en==1'b1)
			r_57_50 <= data_in;
	if (addr_selector[57]&addr_selector[51])
		data_out <= r_57_51;
		if (write_en==1'b1)
			r_57_51 <= data_in;
	if (addr_selector[57]&addr_selector[52])
		data_out <= r_57_52;
		if (write_en==1'b1)
			r_57_52 <= data_in;
	if (addr_selector[57]&addr_selector[53])
		data_out <= r_57_53;
		if (write_en==1'b1)
			r_57_53 <= data_in;
	if (addr_selector[57]&addr_selector[54])
		data_out <= r_57_54;
		if (write_en==1'b1)
			r_57_54 <= data_in;
	if (addr_selector[57]&addr_selector[55])
		data_out <= r_57_55;
		if (write_en==1'b1)
			r_57_55 <= data_in;
	if (addr_selector[57]&addr_selector[56])
		data_out <= r_57_56;
		if (write_en==1'b1)
			r_57_56 <= data_in;
	if (addr_selector[57]&addr_selector[57])
		data_out <= r_57_57;
		if (write_en==1'b1)
			r_57_57 <= data_in;
	if (addr_selector[57]&addr_selector[58])
		data_out <= r_57_58;
		if (write_en==1'b1)
			r_57_58 <= data_in;
	if (addr_selector[57]&addr_selector[59])
		data_out <= r_57_59;
		if (write_en==1'b1)
			r_57_59 <= data_in;
	if (addr_selector[57]&addr_selector[60])
		data_out <= r_57_60;
		if (write_en==1'b1)
			r_57_60 <= data_in;
	if (addr_selector[57]&addr_selector[61])
		data_out <= r_57_61;
		if (write_en==1'b1)
			r_57_61 <= data_in;
	if (addr_selector[57]&addr_selector[62])
		data_out <= r_57_62;
		if (write_en==1'b1)
			r_57_62 <= data_in;
	if (addr_selector[57]&addr_selector[63])
		data_out <= r_57_63;
		if (write_en==1'b1)
			r_57_63 <= data_in;
	if (addr_selector[58]&addr_selector[0])
		data_out <= r_58_0;
		if (write_en==1'b1)
			r_58_0 <= data_in;
	if (addr_selector[58]&addr_selector[1])
		data_out <= r_58_1;
		if (write_en==1'b1)
			r_58_1 <= data_in;
	if (addr_selector[58]&addr_selector[2])
		data_out <= r_58_2;
		if (write_en==1'b1)
			r_58_2 <= data_in;
	if (addr_selector[58]&addr_selector[3])
		data_out <= r_58_3;
		if (write_en==1'b1)
			r_58_3 <= data_in;
	if (addr_selector[58]&addr_selector[4])
		data_out <= r_58_4;
		if (write_en==1'b1)
			r_58_4 <= data_in;
	if (addr_selector[58]&addr_selector[5])
		data_out <= r_58_5;
		if (write_en==1'b1)
			r_58_5 <= data_in;
	if (addr_selector[58]&addr_selector[6])
		data_out <= r_58_6;
		if (write_en==1'b1)
			r_58_6 <= data_in;
	if (addr_selector[58]&addr_selector[7])
		data_out <= r_58_7;
		if (write_en==1'b1)
			r_58_7 <= data_in;
	if (addr_selector[58]&addr_selector[8])
		data_out <= r_58_8;
		if (write_en==1'b1)
			r_58_8 <= data_in;
	if (addr_selector[58]&addr_selector[9])
		data_out <= r_58_9;
		if (write_en==1'b1)
			r_58_9 <= data_in;
	if (addr_selector[58]&addr_selector[10])
		data_out <= r_58_10;
		if (write_en==1'b1)
			r_58_10 <= data_in;
	if (addr_selector[58]&addr_selector[11])
		data_out <= r_58_11;
		if (write_en==1'b1)
			r_58_11 <= data_in;
	if (addr_selector[58]&addr_selector[12])
		data_out <= r_58_12;
		if (write_en==1'b1)
			r_58_12 <= data_in;
	if (addr_selector[58]&addr_selector[13])
		data_out <= r_58_13;
		if (write_en==1'b1)
			r_58_13 <= data_in;
	if (addr_selector[58]&addr_selector[14])
		data_out <= r_58_14;
		if (write_en==1'b1)
			r_58_14 <= data_in;
	if (addr_selector[58]&addr_selector[15])
		data_out <= r_58_15;
		if (write_en==1'b1)
			r_58_15 <= data_in;
	if (addr_selector[58]&addr_selector[16])
		data_out <= r_58_16;
		if (write_en==1'b1)
			r_58_16 <= data_in;
	if (addr_selector[58]&addr_selector[17])
		data_out <= r_58_17;
		if (write_en==1'b1)
			r_58_17 <= data_in;
	if (addr_selector[58]&addr_selector[18])
		data_out <= r_58_18;
		if (write_en==1'b1)
			r_58_18 <= data_in;
	if (addr_selector[58]&addr_selector[19])
		data_out <= r_58_19;
		if (write_en==1'b1)
			r_58_19 <= data_in;
	if (addr_selector[58]&addr_selector[20])
		data_out <= r_58_20;
		if (write_en==1'b1)
			r_58_20 <= data_in;
	if (addr_selector[58]&addr_selector[21])
		data_out <= r_58_21;
		if (write_en==1'b1)
			r_58_21 <= data_in;
	if (addr_selector[58]&addr_selector[22])
		data_out <= r_58_22;
		if (write_en==1'b1)
			r_58_22 <= data_in;
	if (addr_selector[58]&addr_selector[23])
		data_out <= r_58_23;
		if (write_en==1'b1)
			r_58_23 <= data_in;
	if (addr_selector[58]&addr_selector[24])
		data_out <= r_58_24;
		if (write_en==1'b1)
			r_58_24 <= data_in;
	if (addr_selector[58]&addr_selector[25])
		data_out <= r_58_25;
		if (write_en==1'b1)
			r_58_25 <= data_in;
	if (addr_selector[58]&addr_selector[26])
		data_out <= r_58_26;
		if (write_en==1'b1)
			r_58_26 <= data_in;
	if (addr_selector[58]&addr_selector[27])
		data_out <= r_58_27;
		if (write_en==1'b1)
			r_58_27 <= data_in;
	if (addr_selector[58]&addr_selector[28])
		data_out <= r_58_28;
		if (write_en==1'b1)
			r_58_28 <= data_in;
	if (addr_selector[58]&addr_selector[29])
		data_out <= r_58_29;
		if (write_en==1'b1)
			r_58_29 <= data_in;
	if (addr_selector[58]&addr_selector[30])
		data_out <= r_58_30;
		if (write_en==1'b1)
			r_58_30 <= data_in;
	if (addr_selector[58]&addr_selector[31])
		data_out <= r_58_31;
		if (write_en==1'b1)
			r_58_31 <= data_in;
	if (addr_selector[58]&addr_selector[32])
		data_out <= r_58_32;
		if (write_en==1'b1)
			r_58_32 <= data_in;
	if (addr_selector[58]&addr_selector[33])
		data_out <= r_58_33;
		if (write_en==1'b1)
			r_58_33 <= data_in;
	if (addr_selector[58]&addr_selector[34])
		data_out <= r_58_34;
		if (write_en==1'b1)
			r_58_34 <= data_in;
	if (addr_selector[58]&addr_selector[35])
		data_out <= r_58_35;
		if (write_en==1'b1)
			r_58_35 <= data_in;
	if (addr_selector[58]&addr_selector[36])
		data_out <= r_58_36;
		if (write_en==1'b1)
			r_58_36 <= data_in;
	if (addr_selector[58]&addr_selector[37])
		data_out <= r_58_37;
		if (write_en==1'b1)
			r_58_37 <= data_in;
	if (addr_selector[58]&addr_selector[38])
		data_out <= r_58_38;
		if (write_en==1'b1)
			r_58_38 <= data_in;
	if (addr_selector[58]&addr_selector[39])
		data_out <= r_58_39;
		if (write_en==1'b1)
			r_58_39 <= data_in;
	if (addr_selector[58]&addr_selector[40])
		data_out <= r_58_40;
		if (write_en==1'b1)
			r_58_40 <= data_in;
	if (addr_selector[58]&addr_selector[41])
		data_out <= r_58_41;
		if (write_en==1'b1)
			r_58_41 <= data_in;
	if (addr_selector[58]&addr_selector[42])
		data_out <= r_58_42;
		if (write_en==1'b1)
			r_58_42 <= data_in;
	if (addr_selector[58]&addr_selector[43])
		data_out <= r_58_43;
		if (write_en==1'b1)
			r_58_43 <= data_in;
	if (addr_selector[58]&addr_selector[44])
		data_out <= r_58_44;
		if (write_en==1'b1)
			r_58_44 <= data_in;
	if (addr_selector[58]&addr_selector[45])
		data_out <= r_58_45;
		if (write_en==1'b1)
			r_58_45 <= data_in;
	if (addr_selector[58]&addr_selector[46])
		data_out <= r_58_46;
		if (write_en==1'b1)
			r_58_46 <= data_in;
	if (addr_selector[58]&addr_selector[47])
		data_out <= r_58_47;
		if (write_en==1'b1)
			r_58_47 <= data_in;
	if (addr_selector[58]&addr_selector[48])
		data_out <= r_58_48;
		if (write_en==1'b1)
			r_58_48 <= data_in;
	if (addr_selector[58]&addr_selector[49])
		data_out <= r_58_49;
		if (write_en==1'b1)
			r_58_49 <= data_in;
	if (addr_selector[58]&addr_selector[50])
		data_out <= r_58_50;
		if (write_en==1'b1)
			r_58_50 <= data_in;
	if (addr_selector[58]&addr_selector[51])
		data_out <= r_58_51;
		if (write_en==1'b1)
			r_58_51 <= data_in;
	if (addr_selector[58]&addr_selector[52])
		data_out <= r_58_52;
		if (write_en==1'b1)
			r_58_52 <= data_in;
	if (addr_selector[58]&addr_selector[53])
		data_out <= r_58_53;
		if (write_en==1'b1)
			r_58_53 <= data_in;
	if (addr_selector[58]&addr_selector[54])
		data_out <= r_58_54;
		if (write_en==1'b1)
			r_58_54 <= data_in;
	if (addr_selector[58]&addr_selector[55])
		data_out <= r_58_55;
		if (write_en==1'b1)
			r_58_55 <= data_in;
	if (addr_selector[58]&addr_selector[56])
		data_out <= r_58_56;
		if (write_en==1'b1)
			r_58_56 <= data_in;
	if (addr_selector[58]&addr_selector[57])
		data_out <= r_58_57;
		if (write_en==1'b1)
			r_58_57 <= data_in;
	if (addr_selector[58]&addr_selector[58])
		data_out <= r_58_58;
		if (write_en==1'b1)
			r_58_58 <= data_in;
	if (addr_selector[58]&addr_selector[59])
		data_out <= r_58_59;
		if (write_en==1'b1)
			r_58_59 <= data_in;
	if (addr_selector[58]&addr_selector[60])
		data_out <= r_58_60;
		if (write_en==1'b1)
			r_58_60 <= data_in;
	if (addr_selector[58]&addr_selector[61])
		data_out <= r_58_61;
		if (write_en==1'b1)
			r_58_61 <= data_in;
	if (addr_selector[58]&addr_selector[62])
		data_out <= r_58_62;
		if (write_en==1'b1)
			r_58_62 <= data_in;
	if (addr_selector[58]&addr_selector[63])
		data_out <= r_58_63;
		if (write_en==1'b1)
			r_58_63 <= data_in;
	if (addr_selector[59]&addr_selector[0])
		data_out <= r_59_0;
		if (write_en==1'b1)
			r_59_0 <= data_in;
	if (addr_selector[59]&addr_selector[1])
		data_out <= r_59_1;
		if (write_en==1'b1)
			r_59_1 <= data_in;
	if (addr_selector[59]&addr_selector[2])
		data_out <= r_59_2;
		if (write_en==1'b1)
			r_59_2 <= data_in;
	if (addr_selector[59]&addr_selector[3])
		data_out <= r_59_3;
		if (write_en==1'b1)
			r_59_3 <= data_in;
	if (addr_selector[59]&addr_selector[4])
		data_out <= r_59_4;
		if (write_en==1'b1)
			r_59_4 <= data_in;
	if (addr_selector[59]&addr_selector[5])
		data_out <= r_59_5;
		if (write_en==1'b1)
			r_59_5 <= data_in;
	if (addr_selector[59]&addr_selector[6])
		data_out <= r_59_6;
		if (write_en==1'b1)
			r_59_6 <= data_in;
	if (addr_selector[59]&addr_selector[7])
		data_out <= r_59_7;
		if (write_en==1'b1)
			r_59_7 <= data_in;
	if (addr_selector[59]&addr_selector[8])
		data_out <= r_59_8;
		if (write_en==1'b1)
			r_59_8 <= data_in;
	if (addr_selector[59]&addr_selector[9])
		data_out <= r_59_9;
		if (write_en==1'b1)
			r_59_9 <= data_in;
	if (addr_selector[59]&addr_selector[10])
		data_out <= r_59_10;
		if (write_en==1'b1)
			r_59_10 <= data_in;
	if (addr_selector[59]&addr_selector[11])
		data_out <= r_59_11;
		if (write_en==1'b1)
			r_59_11 <= data_in;
	if (addr_selector[59]&addr_selector[12])
		data_out <= r_59_12;
		if (write_en==1'b1)
			r_59_12 <= data_in;
	if (addr_selector[59]&addr_selector[13])
		data_out <= r_59_13;
		if (write_en==1'b1)
			r_59_13 <= data_in;
	if (addr_selector[59]&addr_selector[14])
		data_out <= r_59_14;
		if (write_en==1'b1)
			r_59_14 <= data_in;
	if (addr_selector[59]&addr_selector[15])
		data_out <= r_59_15;
		if (write_en==1'b1)
			r_59_15 <= data_in;
	if (addr_selector[59]&addr_selector[16])
		data_out <= r_59_16;
		if (write_en==1'b1)
			r_59_16 <= data_in;
	if (addr_selector[59]&addr_selector[17])
		data_out <= r_59_17;
		if (write_en==1'b1)
			r_59_17 <= data_in;
	if (addr_selector[59]&addr_selector[18])
		data_out <= r_59_18;
		if (write_en==1'b1)
			r_59_18 <= data_in;
	if (addr_selector[59]&addr_selector[19])
		data_out <= r_59_19;
		if (write_en==1'b1)
			r_59_19 <= data_in;
	if (addr_selector[59]&addr_selector[20])
		data_out <= r_59_20;
		if (write_en==1'b1)
			r_59_20 <= data_in;
	if (addr_selector[59]&addr_selector[21])
		data_out <= r_59_21;
		if (write_en==1'b1)
			r_59_21 <= data_in;
	if (addr_selector[59]&addr_selector[22])
		data_out <= r_59_22;
		if (write_en==1'b1)
			r_59_22 <= data_in;
	if (addr_selector[59]&addr_selector[23])
		data_out <= r_59_23;
		if (write_en==1'b1)
			r_59_23 <= data_in;
	if (addr_selector[59]&addr_selector[24])
		data_out <= r_59_24;
		if (write_en==1'b1)
			r_59_24 <= data_in;
	if (addr_selector[59]&addr_selector[25])
		data_out <= r_59_25;
		if (write_en==1'b1)
			r_59_25 <= data_in;
	if (addr_selector[59]&addr_selector[26])
		data_out <= r_59_26;
		if (write_en==1'b1)
			r_59_26 <= data_in;
	if (addr_selector[59]&addr_selector[27])
		data_out <= r_59_27;
		if (write_en==1'b1)
			r_59_27 <= data_in;
	if (addr_selector[59]&addr_selector[28])
		data_out <= r_59_28;
		if (write_en==1'b1)
			r_59_28 <= data_in;
	if (addr_selector[59]&addr_selector[29])
		data_out <= r_59_29;
		if (write_en==1'b1)
			r_59_29 <= data_in;
	if (addr_selector[59]&addr_selector[30])
		data_out <= r_59_30;
		if (write_en==1'b1)
			r_59_30 <= data_in;
	if (addr_selector[59]&addr_selector[31])
		data_out <= r_59_31;
		if (write_en==1'b1)
			r_59_31 <= data_in;
	if (addr_selector[59]&addr_selector[32])
		data_out <= r_59_32;
		if (write_en==1'b1)
			r_59_32 <= data_in;
	if (addr_selector[59]&addr_selector[33])
		data_out <= r_59_33;
		if (write_en==1'b1)
			r_59_33 <= data_in;
	if (addr_selector[59]&addr_selector[34])
		data_out <= r_59_34;
		if (write_en==1'b1)
			r_59_34 <= data_in;
	if (addr_selector[59]&addr_selector[35])
		data_out <= r_59_35;
		if (write_en==1'b1)
			r_59_35 <= data_in;
	if (addr_selector[59]&addr_selector[36])
		data_out <= r_59_36;
		if (write_en==1'b1)
			r_59_36 <= data_in;
	if (addr_selector[59]&addr_selector[37])
		data_out <= r_59_37;
		if (write_en==1'b1)
			r_59_37 <= data_in;
	if (addr_selector[59]&addr_selector[38])
		data_out <= r_59_38;
		if (write_en==1'b1)
			r_59_38 <= data_in;
	if (addr_selector[59]&addr_selector[39])
		data_out <= r_59_39;
		if (write_en==1'b1)
			r_59_39 <= data_in;
	if (addr_selector[59]&addr_selector[40])
		data_out <= r_59_40;
		if (write_en==1'b1)
			r_59_40 <= data_in;
	if (addr_selector[59]&addr_selector[41])
		data_out <= r_59_41;
		if (write_en==1'b1)
			r_59_41 <= data_in;
	if (addr_selector[59]&addr_selector[42])
		data_out <= r_59_42;
		if (write_en==1'b1)
			r_59_42 <= data_in;
	if (addr_selector[59]&addr_selector[43])
		data_out <= r_59_43;
		if (write_en==1'b1)
			r_59_43 <= data_in;
	if (addr_selector[59]&addr_selector[44])
		data_out <= r_59_44;
		if (write_en==1'b1)
			r_59_44 <= data_in;
	if (addr_selector[59]&addr_selector[45])
		data_out <= r_59_45;
		if (write_en==1'b1)
			r_59_45 <= data_in;
	if (addr_selector[59]&addr_selector[46])
		data_out <= r_59_46;
		if (write_en==1'b1)
			r_59_46 <= data_in;
	if (addr_selector[59]&addr_selector[47])
		data_out <= r_59_47;
		if (write_en==1'b1)
			r_59_47 <= data_in;
	if (addr_selector[59]&addr_selector[48])
		data_out <= r_59_48;
		if (write_en==1'b1)
			r_59_48 <= data_in;
	if (addr_selector[59]&addr_selector[49])
		data_out <= r_59_49;
		if (write_en==1'b1)
			r_59_49 <= data_in;
	if (addr_selector[59]&addr_selector[50])
		data_out <= r_59_50;
		if (write_en==1'b1)
			r_59_50 <= data_in;
	if (addr_selector[59]&addr_selector[51])
		data_out <= r_59_51;
		if (write_en==1'b1)
			r_59_51 <= data_in;
	if (addr_selector[59]&addr_selector[52])
		data_out <= r_59_52;
		if (write_en==1'b1)
			r_59_52 <= data_in;
	if (addr_selector[59]&addr_selector[53])
		data_out <= r_59_53;
		if (write_en==1'b1)
			r_59_53 <= data_in;
	if (addr_selector[59]&addr_selector[54])
		data_out <= r_59_54;
		if (write_en==1'b1)
			r_59_54 <= data_in;
	if (addr_selector[59]&addr_selector[55])
		data_out <= r_59_55;
		if (write_en==1'b1)
			r_59_55 <= data_in;
	if (addr_selector[59]&addr_selector[56])
		data_out <= r_59_56;
		if (write_en==1'b1)
			r_59_56 <= data_in;
	if (addr_selector[59]&addr_selector[57])
		data_out <= r_59_57;
		if (write_en==1'b1)
			r_59_57 <= data_in;
	if (addr_selector[59]&addr_selector[58])
		data_out <= r_59_58;
		if (write_en==1'b1)
			r_59_58 <= data_in;
	if (addr_selector[59]&addr_selector[59])
		data_out <= r_59_59;
		if (write_en==1'b1)
			r_59_59 <= data_in;
	if (addr_selector[59]&addr_selector[60])
		data_out <= r_59_60;
		if (write_en==1'b1)
			r_59_60 <= data_in;
	if (addr_selector[59]&addr_selector[61])
		data_out <= r_59_61;
		if (write_en==1'b1)
			r_59_61 <= data_in;
	if (addr_selector[59]&addr_selector[62])
		data_out <= r_59_62;
		if (write_en==1'b1)
			r_59_62 <= data_in;
	if (addr_selector[59]&addr_selector[63])
		data_out <= r_59_63;
		if (write_en==1'b1)
			r_59_63 <= data_in;
	if (addr_selector[60]&addr_selector[0])
		data_out <= r_60_0;
		if (write_en==1'b1)
			r_60_0 <= data_in;
	if (addr_selector[60]&addr_selector[1])
		data_out <= r_60_1;
		if (write_en==1'b1)
			r_60_1 <= data_in;
	if (addr_selector[60]&addr_selector[2])
		data_out <= r_60_2;
		if (write_en==1'b1)
			r_60_2 <= data_in;
	if (addr_selector[60]&addr_selector[3])
		data_out <= r_60_3;
		if (write_en==1'b1)
			r_60_3 <= data_in;
	if (addr_selector[60]&addr_selector[4])
		data_out <= r_60_4;
		if (write_en==1'b1)
			r_60_4 <= data_in;
	if (addr_selector[60]&addr_selector[5])
		data_out <= r_60_5;
		if (write_en==1'b1)
			r_60_5 <= data_in;
	if (addr_selector[60]&addr_selector[6])
		data_out <= r_60_6;
		if (write_en==1'b1)
			r_60_6 <= data_in;
	if (addr_selector[60]&addr_selector[7])
		data_out <= r_60_7;
		if (write_en==1'b1)
			r_60_7 <= data_in;
	if (addr_selector[60]&addr_selector[8])
		data_out <= r_60_8;
		if (write_en==1'b1)
			r_60_8 <= data_in;
	if (addr_selector[60]&addr_selector[9])
		data_out <= r_60_9;
		if (write_en==1'b1)
			r_60_9 <= data_in;
	if (addr_selector[60]&addr_selector[10])
		data_out <= r_60_10;
		if (write_en==1'b1)
			r_60_10 <= data_in;
	if (addr_selector[60]&addr_selector[11])
		data_out <= r_60_11;
		if (write_en==1'b1)
			r_60_11 <= data_in;
	if (addr_selector[60]&addr_selector[12])
		data_out <= r_60_12;
		if (write_en==1'b1)
			r_60_12 <= data_in;
	if (addr_selector[60]&addr_selector[13])
		data_out <= r_60_13;
		if (write_en==1'b1)
			r_60_13 <= data_in;
	if (addr_selector[60]&addr_selector[14])
		data_out <= r_60_14;
		if (write_en==1'b1)
			r_60_14 <= data_in;
	if (addr_selector[60]&addr_selector[15])
		data_out <= r_60_15;
		if (write_en==1'b1)
			r_60_15 <= data_in;
	if (addr_selector[60]&addr_selector[16])
		data_out <= r_60_16;
		if (write_en==1'b1)
			r_60_16 <= data_in;
	if (addr_selector[60]&addr_selector[17])
		data_out <= r_60_17;
		if (write_en==1'b1)
			r_60_17 <= data_in;
	if (addr_selector[60]&addr_selector[18])
		data_out <= r_60_18;
		if (write_en==1'b1)
			r_60_18 <= data_in;
	if (addr_selector[60]&addr_selector[19])
		data_out <= r_60_19;
		if (write_en==1'b1)
			r_60_19 <= data_in;
	if (addr_selector[60]&addr_selector[20])
		data_out <= r_60_20;
		if (write_en==1'b1)
			r_60_20 <= data_in;
	if (addr_selector[60]&addr_selector[21])
		data_out <= r_60_21;
		if (write_en==1'b1)
			r_60_21 <= data_in;
	if (addr_selector[60]&addr_selector[22])
		data_out <= r_60_22;
		if (write_en==1'b1)
			r_60_22 <= data_in;
	if (addr_selector[60]&addr_selector[23])
		data_out <= r_60_23;
		if (write_en==1'b1)
			r_60_23 <= data_in;
	if (addr_selector[60]&addr_selector[24])
		data_out <= r_60_24;
		if (write_en==1'b1)
			r_60_24 <= data_in;
	if (addr_selector[60]&addr_selector[25])
		data_out <= r_60_25;
		if (write_en==1'b1)
			r_60_25 <= data_in;
	if (addr_selector[60]&addr_selector[26])
		data_out <= r_60_26;
		if (write_en==1'b1)
			r_60_26 <= data_in;
	if (addr_selector[60]&addr_selector[27])
		data_out <= r_60_27;
		if (write_en==1'b1)
			r_60_27 <= data_in;
	if (addr_selector[60]&addr_selector[28])
		data_out <= r_60_28;
		if (write_en==1'b1)
			r_60_28 <= data_in;
	if (addr_selector[60]&addr_selector[29])
		data_out <= r_60_29;
		if (write_en==1'b1)
			r_60_29 <= data_in;
	if (addr_selector[60]&addr_selector[30])
		data_out <= r_60_30;
		if (write_en==1'b1)
			r_60_30 <= data_in;
	if (addr_selector[60]&addr_selector[31])
		data_out <= r_60_31;
		if (write_en==1'b1)
			r_60_31 <= data_in;
	if (addr_selector[60]&addr_selector[32])
		data_out <= r_60_32;
		if (write_en==1'b1)
			r_60_32 <= data_in;
	if (addr_selector[60]&addr_selector[33])
		data_out <= r_60_33;
		if (write_en==1'b1)
			r_60_33 <= data_in;
	if (addr_selector[60]&addr_selector[34])
		data_out <= r_60_34;
		if (write_en==1'b1)
			r_60_34 <= data_in;
	if (addr_selector[60]&addr_selector[35])
		data_out <= r_60_35;
		if (write_en==1'b1)
			r_60_35 <= data_in;
	if (addr_selector[60]&addr_selector[36])
		data_out <= r_60_36;
		if (write_en==1'b1)
			r_60_36 <= data_in;
	if (addr_selector[60]&addr_selector[37])
		data_out <= r_60_37;
		if (write_en==1'b1)
			r_60_37 <= data_in;
	if (addr_selector[60]&addr_selector[38])
		data_out <= r_60_38;
		if (write_en==1'b1)
			r_60_38 <= data_in;
	if (addr_selector[60]&addr_selector[39])
		data_out <= r_60_39;
		if (write_en==1'b1)
			r_60_39 <= data_in;
	if (addr_selector[60]&addr_selector[40])
		data_out <= r_60_40;
		if (write_en==1'b1)
			r_60_40 <= data_in;
	if (addr_selector[60]&addr_selector[41])
		data_out <= r_60_41;
		if (write_en==1'b1)
			r_60_41 <= data_in;
	if (addr_selector[60]&addr_selector[42])
		data_out <= r_60_42;
		if (write_en==1'b1)
			r_60_42 <= data_in;
	if (addr_selector[60]&addr_selector[43])
		data_out <= r_60_43;
		if (write_en==1'b1)
			r_60_43 <= data_in;
	if (addr_selector[60]&addr_selector[44])
		data_out <= r_60_44;
		if (write_en==1'b1)
			r_60_44 <= data_in;
	if (addr_selector[60]&addr_selector[45])
		data_out <= r_60_45;
		if (write_en==1'b1)
			r_60_45 <= data_in;
	if (addr_selector[60]&addr_selector[46])
		data_out <= r_60_46;
		if (write_en==1'b1)
			r_60_46 <= data_in;
	if (addr_selector[60]&addr_selector[47])
		data_out <= r_60_47;
		if (write_en==1'b1)
			r_60_47 <= data_in;
	if (addr_selector[60]&addr_selector[48])
		data_out <= r_60_48;
		if (write_en==1'b1)
			r_60_48 <= data_in;
	if (addr_selector[60]&addr_selector[49])
		data_out <= r_60_49;
		if (write_en==1'b1)
			r_60_49 <= data_in;
	if (addr_selector[60]&addr_selector[50])
		data_out <= r_60_50;
		if (write_en==1'b1)
			r_60_50 <= data_in;
	if (addr_selector[60]&addr_selector[51])
		data_out <= r_60_51;
		if (write_en==1'b1)
			r_60_51 <= data_in;
	if (addr_selector[60]&addr_selector[52])
		data_out <= r_60_52;
		if (write_en==1'b1)
			r_60_52 <= data_in;
	if (addr_selector[60]&addr_selector[53])
		data_out <= r_60_53;
		if (write_en==1'b1)
			r_60_53 <= data_in;
	if (addr_selector[60]&addr_selector[54])
		data_out <= r_60_54;
		if (write_en==1'b1)
			r_60_54 <= data_in;
	if (addr_selector[60]&addr_selector[55])
		data_out <= r_60_55;
		if (write_en==1'b1)
			r_60_55 <= data_in;
	if (addr_selector[60]&addr_selector[56])
		data_out <= r_60_56;
		if (write_en==1'b1)
			r_60_56 <= data_in;
	if (addr_selector[60]&addr_selector[57])
		data_out <= r_60_57;
		if (write_en==1'b1)
			r_60_57 <= data_in;
	if (addr_selector[60]&addr_selector[58])
		data_out <= r_60_58;
		if (write_en==1'b1)
			r_60_58 <= data_in;
	if (addr_selector[60]&addr_selector[59])
		data_out <= r_60_59;
		if (write_en==1'b1)
			r_60_59 <= data_in;
	if (addr_selector[60]&addr_selector[60])
		data_out <= r_60_60;
		if (write_en==1'b1)
			r_60_60 <= data_in;
	if (addr_selector[60]&addr_selector[61])
		data_out <= r_60_61;
		if (write_en==1'b1)
			r_60_61 <= data_in;
	if (addr_selector[60]&addr_selector[62])
		data_out <= r_60_62;
		if (write_en==1'b1)
			r_60_62 <= data_in;
	if (addr_selector[60]&addr_selector[63])
		data_out <= r_60_63;
		if (write_en==1'b1)
			r_60_63 <= data_in;
	if (addr_selector[61]&addr_selector[0])
		data_out <= r_61_0;
		if (write_en==1'b1)
			r_61_0 <= data_in;
	if (addr_selector[61]&addr_selector[1])
		data_out <= r_61_1;
		if (write_en==1'b1)
			r_61_1 <= data_in;
	if (addr_selector[61]&addr_selector[2])
		data_out <= r_61_2;
		if (write_en==1'b1)
			r_61_2 <= data_in;
	if (addr_selector[61]&addr_selector[3])
		data_out <= r_61_3;
		if (write_en==1'b1)
			r_61_3 <= data_in;
	if (addr_selector[61]&addr_selector[4])
		data_out <= r_61_4;
		if (write_en==1'b1)
			r_61_4 <= data_in;
	if (addr_selector[61]&addr_selector[5])
		data_out <= r_61_5;
		if (write_en==1'b1)
			r_61_5 <= data_in;
	if (addr_selector[61]&addr_selector[6])
		data_out <= r_61_6;
		if (write_en==1'b1)
			r_61_6 <= data_in;
	if (addr_selector[61]&addr_selector[7])
		data_out <= r_61_7;
		if (write_en==1'b1)
			r_61_7 <= data_in;
	if (addr_selector[61]&addr_selector[8])
		data_out <= r_61_8;
		if (write_en==1'b1)
			r_61_8 <= data_in;
	if (addr_selector[61]&addr_selector[9])
		data_out <= r_61_9;
		if (write_en==1'b1)
			r_61_9 <= data_in;
	if (addr_selector[61]&addr_selector[10])
		data_out <= r_61_10;
		if (write_en==1'b1)
			r_61_10 <= data_in;
	if (addr_selector[61]&addr_selector[11])
		data_out <= r_61_11;
		if (write_en==1'b1)
			r_61_11 <= data_in;
	if (addr_selector[61]&addr_selector[12])
		data_out <= r_61_12;
		if (write_en==1'b1)
			r_61_12 <= data_in;
	if (addr_selector[61]&addr_selector[13])
		data_out <= r_61_13;
		if (write_en==1'b1)
			r_61_13 <= data_in;
	if (addr_selector[61]&addr_selector[14])
		data_out <= r_61_14;
		if (write_en==1'b1)
			r_61_14 <= data_in;
	if (addr_selector[61]&addr_selector[15])
		data_out <= r_61_15;
		if (write_en==1'b1)
			r_61_15 <= data_in;
	if (addr_selector[61]&addr_selector[16])
		data_out <= r_61_16;
		if (write_en==1'b1)
			r_61_16 <= data_in;
	if (addr_selector[61]&addr_selector[17])
		data_out <= r_61_17;
		if (write_en==1'b1)
			r_61_17 <= data_in;
	if (addr_selector[61]&addr_selector[18])
		data_out <= r_61_18;
		if (write_en==1'b1)
			r_61_18 <= data_in;
	if (addr_selector[61]&addr_selector[19])
		data_out <= r_61_19;
		if (write_en==1'b1)
			r_61_19 <= data_in;
	if (addr_selector[61]&addr_selector[20])
		data_out <= r_61_20;
		if (write_en==1'b1)
			r_61_20 <= data_in;
	if (addr_selector[61]&addr_selector[21])
		data_out <= r_61_21;
		if (write_en==1'b1)
			r_61_21 <= data_in;
	if (addr_selector[61]&addr_selector[22])
		data_out <= r_61_22;
		if (write_en==1'b1)
			r_61_22 <= data_in;
	if (addr_selector[61]&addr_selector[23])
		data_out <= r_61_23;
		if (write_en==1'b1)
			r_61_23 <= data_in;
	if (addr_selector[61]&addr_selector[24])
		data_out <= r_61_24;
		if (write_en==1'b1)
			r_61_24 <= data_in;
	if (addr_selector[61]&addr_selector[25])
		data_out <= r_61_25;
		if (write_en==1'b1)
			r_61_25 <= data_in;
	if (addr_selector[61]&addr_selector[26])
		data_out <= r_61_26;
		if (write_en==1'b1)
			r_61_26 <= data_in;
	if (addr_selector[61]&addr_selector[27])
		data_out <= r_61_27;
		if (write_en==1'b1)
			r_61_27 <= data_in;
	if (addr_selector[61]&addr_selector[28])
		data_out <= r_61_28;
		if (write_en==1'b1)
			r_61_28 <= data_in;
	if (addr_selector[61]&addr_selector[29])
		data_out <= r_61_29;
		if (write_en==1'b1)
			r_61_29 <= data_in;
	if (addr_selector[61]&addr_selector[30])
		data_out <= r_61_30;
		if (write_en==1'b1)
			r_61_30 <= data_in;
	if (addr_selector[61]&addr_selector[31])
		data_out <= r_61_31;
		if (write_en==1'b1)
			r_61_31 <= data_in;
	if (addr_selector[61]&addr_selector[32])
		data_out <= r_61_32;
		if (write_en==1'b1)
			r_61_32 <= data_in;
	if (addr_selector[61]&addr_selector[33])
		data_out <= r_61_33;
		if (write_en==1'b1)
			r_61_33 <= data_in;
	if (addr_selector[61]&addr_selector[34])
		data_out <= r_61_34;
		if (write_en==1'b1)
			r_61_34 <= data_in;
	if (addr_selector[61]&addr_selector[35])
		data_out <= r_61_35;
		if (write_en==1'b1)
			r_61_35 <= data_in;
	if (addr_selector[61]&addr_selector[36])
		data_out <= r_61_36;
		if (write_en==1'b1)
			r_61_36 <= data_in;
	if (addr_selector[61]&addr_selector[37])
		data_out <= r_61_37;
		if (write_en==1'b1)
			r_61_37 <= data_in;
	if (addr_selector[61]&addr_selector[38])
		data_out <= r_61_38;
		if (write_en==1'b1)
			r_61_38 <= data_in;
	if (addr_selector[61]&addr_selector[39])
		data_out <= r_61_39;
		if (write_en==1'b1)
			r_61_39 <= data_in;
	if (addr_selector[61]&addr_selector[40])
		data_out <= r_61_40;
		if (write_en==1'b1)
			r_61_40 <= data_in;
	if (addr_selector[61]&addr_selector[41])
		data_out <= r_61_41;
		if (write_en==1'b1)
			r_61_41 <= data_in;
	if (addr_selector[61]&addr_selector[42])
		data_out <= r_61_42;
		if (write_en==1'b1)
			r_61_42 <= data_in;
	if (addr_selector[61]&addr_selector[43])
		data_out <= r_61_43;
		if (write_en==1'b1)
			r_61_43 <= data_in;
	if (addr_selector[61]&addr_selector[44])
		data_out <= r_61_44;
		if (write_en==1'b1)
			r_61_44 <= data_in;
	if (addr_selector[61]&addr_selector[45])
		data_out <= r_61_45;
		if (write_en==1'b1)
			r_61_45 <= data_in;
	if (addr_selector[61]&addr_selector[46])
		data_out <= r_61_46;
		if (write_en==1'b1)
			r_61_46 <= data_in;
	if (addr_selector[61]&addr_selector[47])
		data_out <= r_61_47;
		if (write_en==1'b1)
			r_61_47 <= data_in;
	if (addr_selector[61]&addr_selector[48])
		data_out <= r_61_48;
		if (write_en==1'b1)
			r_61_48 <= data_in;
	if (addr_selector[61]&addr_selector[49])
		data_out <= r_61_49;
		if (write_en==1'b1)
			r_61_49 <= data_in;
	if (addr_selector[61]&addr_selector[50])
		data_out <= r_61_50;
		if (write_en==1'b1)
			r_61_50 <= data_in;
	if (addr_selector[61]&addr_selector[51])
		data_out <= r_61_51;
		if (write_en==1'b1)
			r_61_51 <= data_in;
	if (addr_selector[61]&addr_selector[52])
		data_out <= r_61_52;
		if (write_en==1'b1)
			r_61_52 <= data_in;
	if (addr_selector[61]&addr_selector[53])
		data_out <= r_61_53;
		if (write_en==1'b1)
			r_61_53 <= data_in;
	if (addr_selector[61]&addr_selector[54])
		data_out <= r_61_54;
		if (write_en==1'b1)
			r_61_54 <= data_in;
	if (addr_selector[61]&addr_selector[55])
		data_out <= r_61_55;
		if (write_en==1'b1)
			r_61_55 <= data_in;
	if (addr_selector[61]&addr_selector[56])
		data_out <= r_61_56;
		if (write_en==1'b1)
			r_61_56 <= data_in;
	if (addr_selector[61]&addr_selector[57])
		data_out <= r_61_57;
		if (write_en==1'b1)
			r_61_57 <= data_in;
	if (addr_selector[61]&addr_selector[58])
		data_out <= r_61_58;
		if (write_en==1'b1)
			r_61_58 <= data_in;
	if (addr_selector[61]&addr_selector[59])
		data_out <= r_61_59;
		if (write_en==1'b1)
			r_61_59 <= data_in;
	if (addr_selector[61]&addr_selector[60])
		data_out <= r_61_60;
		if (write_en==1'b1)
			r_61_60 <= data_in;
	if (addr_selector[61]&addr_selector[61])
		data_out <= r_61_61;
		if (write_en==1'b1)
			r_61_61 <= data_in;
	if (addr_selector[61]&addr_selector[62])
		data_out <= r_61_62;
		if (write_en==1'b1)
			r_61_62 <= data_in;
	if (addr_selector[61]&addr_selector[63])
		data_out <= r_61_63;
		if (write_en==1'b1)
			r_61_63 <= data_in;
	if (addr_selector[62]&addr_selector[0])
		data_out <= r_62_0;
		if (write_en==1'b1)
			r_62_0 <= data_in;
	if (addr_selector[62]&addr_selector[1])
		data_out <= r_62_1;
		if (write_en==1'b1)
			r_62_1 <= data_in;
	if (addr_selector[62]&addr_selector[2])
		data_out <= r_62_2;
		if (write_en==1'b1)
			r_62_2 <= data_in;
	if (addr_selector[62]&addr_selector[3])
		data_out <= r_62_3;
		if (write_en==1'b1)
			r_62_3 <= data_in;
	if (addr_selector[62]&addr_selector[4])
		data_out <= r_62_4;
		if (write_en==1'b1)
			r_62_4 <= data_in;
	if (addr_selector[62]&addr_selector[5])
		data_out <= r_62_5;
		if (write_en==1'b1)
			r_62_5 <= data_in;
	if (addr_selector[62]&addr_selector[6])
		data_out <= r_62_6;
		if (write_en==1'b1)
			r_62_6 <= data_in;
	if (addr_selector[62]&addr_selector[7])
		data_out <= r_62_7;
		if (write_en==1'b1)
			r_62_7 <= data_in;
	if (addr_selector[62]&addr_selector[8])
		data_out <= r_62_8;
		if (write_en==1'b1)
			r_62_8 <= data_in;
	if (addr_selector[62]&addr_selector[9])
		data_out <= r_62_9;
		if (write_en==1'b1)
			r_62_9 <= data_in;
	if (addr_selector[62]&addr_selector[10])
		data_out <= r_62_10;
		if (write_en==1'b1)
			r_62_10 <= data_in;
	if (addr_selector[62]&addr_selector[11])
		data_out <= r_62_11;
		if (write_en==1'b1)
			r_62_11 <= data_in;
	if (addr_selector[62]&addr_selector[12])
		data_out <= r_62_12;
		if (write_en==1'b1)
			r_62_12 <= data_in;
	if (addr_selector[62]&addr_selector[13])
		data_out <= r_62_13;
		if (write_en==1'b1)
			r_62_13 <= data_in;
	if (addr_selector[62]&addr_selector[14])
		data_out <= r_62_14;
		if (write_en==1'b1)
			r_62_14 <= data_in;
	if (addr_selector[62]&addr_selector[15])
		data_out <= r_62_15;
		if (write_en==1'b1)
			r_62_15 <= data_in;
	if (addr_selector[62]&addr_selector[16])
		data_out <= r_62_16;
		if (write_en==1'b1)
			r_62_16 <= data_in;
	if (addr_selector[62]&addr_selector[17])
		data_out <= r_62_17;
		if (write_en==1'b1)
			r_62_17 <= data_in;
	if (addr_selector[62]&addr_selector[18])
		data_out <= r_62_18;
		if (write_en==1'b1)
			r_62_18 <= data_in;
	if (addr_selector[62]&addr_selector[19])
		data_out <= r_62_19;
		if (write_en==1'b1)
			r_62_19 <= data_in;
	if (addr_selector[62]&addr_selector[20])
		data_out <= r_62_20;
		if (write_en==1'b1)
			r_62_20 <= data_in;
	if (addr_selector[62]&addr_selector[21])
		data_out <= r_62_21;
		if (write_en==1'b1)
			r_62_21 <= data_in;
	if (addr_selector[62]&addr_selector[22])
		data_out <= r_62_22;
		if (write_en==1'b1)
			r_62_22 <= data_in;
	if (addr_selector[62]&addr_selector[23])
		data_out <= r_62_23;
		if (write_en==1'b1)
			r_62_23 <= data_in;
	if (addr_selector[62]&addr_selector[24])
		data_out <= r_62_24;
		if (write_en==1'b1)
			r_62_24 <= data_in;
	if (addr_selector[62]&addr_selector[25])
		data_out <= r_62_25;
		if (write_en==1'b1)
			r_62_25 <= data_in;
	if (addr_selector[62]&addr_selector[26])
		data_out <= r_62_26;
		if (write_en==1'b1)
			r_62_26 <= data_in;
	if (addr_selector[62]&addr_selector[27])
		data_out <= r_62_27;
		if (write_en==1'b1)
			r_62_27 <= data_in;
	if (addr_selector[62]&addr_selector[28])
		data_out <= r_62_28;
		if (write_en==1'b1)
			r_62_28 <= data_in;
	if (addr_selector[62]&addr_selector[29])
		data_out <= r_62_29;
		if (write_en==1'b1)
			r_62_29 <= data_in;
	if (addr_selector[62]&addr_selector[30])
		data_out <= r_62_30;
		if (write_en==1'b1)
			r_62_30 <= data_in;
	if (addr_selector[62]&addr_selector[31])
		data_out <= r_62_31;
		if (write_en==1'b1)
			r_62_31 <= data_in;
	if (addr_selector[62]&addr_selector[32])
		data_out <= r_62_32;
		if (write_en==1'b1)
			r_62_32 <= data_in;
	if (addr_selector[62]&addr_selector[33])
		data_out <= r_62_33;
		if (write_en==1'b1)
			r_62_33 <= data_in;
	if (addr_selector[62]&addr_selector[34])
		data_out <= r_62_34;
		if (write_en==1'b1)
			r_62_34 <= data_in;
	if (addr_selector[62]&addr_selector[35])
		data_out <= r_62_35;
		if (write_en==1'b1)
			r_62_35 <= data_in;
	if (addr_selector[62]&addr_selector[36])
		data_out <= r_62_36;
		if (write_en==1'b1)
			r_62_36 <= data_in;
	if (addr_selector[62]&addr_selector[37])
		data_out <= r_62_37;
		if (write_en==1'b1)
			r_62_37 <= data_in;
	if (addr_selector[62]&addr_selector[38])
		data_out <= r_62_38;
		if (write_en==1'b1)
			r_62_38 <= data_in;
	if (addr_selector[62]&addr_selector[39])
		data_out <= r_62_39;
		if (write_en==1'b1)
			r_62_39 <= data_in;
	if (addr_selector[62]&addr_selector[40])
		data_out <= r_62_40;
		if (write_en==1'b1)
			r_62_40 <= data_in;
	if (addr_selector[62]&addr_selector[41])
		data_out <= r_62_41;
		if (write_en==1'b1)
			r_62_41 <= data_in;
	if (addr_selector[62]&addr_selector[42])
		data_out <= r_62_42;
		if (write_en==1'b1)
			r_62_42 <= data_in;
	if (addr_selector[62]&addr_selector[43])
		data_out <= r_62_43;
		if (write_en==1'b1)
			r_62_43 <= data_in;
	if (addr_selector[62]&addr_selector[44])
		data_out <= r_62_44;
		if (write_en==1'b1)
			r_62_44 <= data_in;
	if (addr_selector[62]&addr_selector[45])
		data_out <= r_62_45;
		if (write_en==1'b1)
			r_62_45 <= data_in;
	if (addr_selector[62]&addr_selector[46])
		data_out <= r_62_46;
		if (write_en==1'b1)
			r_62_46 <= data_in;
	if (addr_selector[62]&addr_selector[47])
		data_out <= r_62_47;
		if (write_en==1'b1)
			r_62_47 <= data_in;
	if (addr_selector[62]&addr_selector[48])
		data_out <= r_62_48;
		if (write_en==1'b1)
			r_62_48 <= data_in;
	if (addr_selector[62]&addr_selector[49])
		data_out <= r_62_49;
		if (write_en==1'b1)
			r_62_49 <= data_in;
	if (addr_selector[62]&addr_selector[50])
		data_out <= r_62_50;
		if (write_en==1'b1)
			r_62_50 <= data_in;
	if (addr_selector[62]&addr_selector[51])
		data_out <= r_62_51;
		if (write_en==1'b1)
			r_62_51 <= data_in;
	if (addr_selector[62]&addr_selector[52])
		data_out <= r_62_52;
		if (write_en==1'b1)
			r_62_52 <= data_in;
	if (addr_selector[62]&addr_selector[53])
		data_out <= r_62_53;
		if (write_en==1'b1)
			r_62_53 <= data_in;
	if (addr_selector[62]&addr_selector[54])
		data_out <= r_62_54;
		if (write_en==1'b1)
			r_62_54 <= data_in;
	if (addr_selector[62]&addr_selector[55])
		data_out <= r_62_55;
		if (write_en==1'b1)
			r_62_55 <= data_in;
	if (addr_selector[62]&addr_selector[56])
		data_out <= r_62_56;
		if (write_en==1'b1)
			r_62_56 <= data_in;
	if (addr_selector[62]&addr_selector[57])
		data_out <= r_62_57;
		if (write_en==1'b1)
			r_62_57 <= data_in;
	if (addr_selector[62]&addr_selector[58])
		data_out <= r_62_58;
		if (write_en==1'b1)
			r_62_58 <= data_in;
	if (addr_selector[62]&addr_selector[59])
		data_out <= r_62_59;
		if (write_en==1'b1)
			r_62_59 <= data_in;
	if (addr_selector[62]&addr_selector[60])
		data_out <= r_62_60;
		if (write_en==1'b1)
			r_62_60 <= data_in;
	if (addr_selector[62]&addr_selector[61])
		data_out <= r_62_61;
		if (write_en==1'b1)
			r_62_61 <= data_in;
	if (addr_selector[62]&addr_selector[62])
		data_out <= r_62_62;
		if (write_en==1'b1)
			r_62_62 <= data_in;
	if (addr_selector[62]&addr_selector[63])
		data_out <= r_62_63;
		if (write_en==1'b1)
			r_62_63 <= data_in;
	if (addr_selector[63]&addr_selector[0])
		data_out <= r_63_0;
		if (write_en==1'b1)
			r_63_0 <= data_in;
	if (addr_selector[63]&addr_selector[1])
		data_out <= r_63_1;
		if (write_en==1'b1)
			r_63_1 <= data_in;
	if (addr_selector[63]&addr_selector[2])
		data_out <= r_63_2;
		if (write_en==1'b1)
			r_63_2 <= data_in;
	if (addr_selector[63]&addr_selector[3])
		data_out <= r_63_3;
		if (write_en==1'b1)
			r_63_3 <= data_in;
	if (addr_selector[63]&addr_selector[4])
		data_out <= r_63_4;
		if (write_en==1'b1)
			r_63_4 <= data_in;
	if (addr_selector[63]&addr_selector[5])
		data_out <= r_63_5;
		if (write_en==1'b1)
			r_63_5 <= data_in;
	if (addr_selector[63]&addr_selector[6])
		data_out <= r_63_6;
		if (write_en==1'b1)
			r_63_6 <= data_in;
	if (addr_selector[63]&addr_selector[7])
		data_out <= r_63_7;
		if (write_en==1'b1)
			r_63_7 <= data_in;
	if (addr_selector[63]&addr_selector[8])
		data_out <= r_63_8;
		if (write_en==1'b1)
			r_63_8 <= data_in;
	if (addr_selector[63]&addr_selector[9])
		data_out <= r_63_9;
		if (write_en==1'b1)
			r_63_9 <= data_in;
	if (addr_selector[63]&addr_selector[10])
		data_out <= r_63_10;
		if (write_en==1'b1)
			r_63_10 <= data_in;
	if (addr_selector[63]&addr_selector[11])
		data_out <= r_63_11;
		if (write_en==1'b1)
			r_63_11 <= data_in;
	if (addr_selector[63]&addr_selector[12])
		data_out <= r_63_12;
		if (write_en==1'b1)
			r_63_12 <= data_in;
	if (addr_selector[63]&addr_selector[13])
		data_out <= r_63_13;
		if (write_en==1'b1)
			r_63_13 <= data_in;
	if (addr_selector[63]&addr_selector[14])
		data_out <= r_63_14;
		if (write_en==1'b1)
			r_63_14 <= data_in;
	if (addr_selector[63]&addr_selector[15])
		data_out <= r_63_15;
		if (write_en==1'b1)
			r_63_15 <= data_in;
	if (addr_selector[63]&addr_selector[16])
		data_out <= r_63_16;
		if (write_en==1'b1)
			r_63_16 <= data_in;
	if (addr_selector[63]&addr_selector[17])
		data_out <= r_63_17;
		if (write_en==1'b1)
			r_63_17 <= data_in;
	if (addr_selector[63]&addr_selector[18])
		data_out <= r_63_18;
		if (write_en==1'b1)
			r_63_18 <= data_in;
	if (addr_selector[63]&addr_selector[19])
		data_out <= r_63_19;
		if (write_en==1'b1)
			r_63_19 <= data_in;
	if (addr_selector[63]&addr_selector[20])
		data_out <= r_63_20;
		if (write_en==1'b1)
			r_63_20 <= data_in;
	if (addr_selector[63]&addr_selector[21])
		data_out <= r_63_21;
		if (write_en==1'b1)
			r_63_21 <= data_in;
	if (addr_selector[63]&addr_selector[22])
		data_out <= r_63_22;
		if (write_en==1'b1)
			r_63_22 <= data_in;
	if (addr_selector[63]&addr_selector[23])
		data_out <= r_63_23;
		if (write_en==1'b1)
			r_63_23 <= data_in;
	if (addr_selector[63]&addr_selector[24])
		data_out <= r_63_24;
		if (write_en==1'b1)
			r_63_24 <= data_in;
	if (addr_selector[63]&addr_selector[25])
		data_out <= r_63_25;
		if (write_en==1'b1)
			r_63_25 <= data_in;
	if (addr_selector[63]&addr_selector[26])
		data_out <= r_63_26;
		if (write_en==1'b1)
			r_63_26 <= data_in;
	if (addr_selector[63]&addr_selector[27])
		data_out <= r_63_27;
		if (write_en==1'b1)
			r_63_27 <= data_in;
	if (addr_selector[63]&addr_selector[28])
		data_out <= r_63_28;
		if (write_en==1'b1)
			r_63_28 <= data_in;
	if (addr_selector[63]&addr_selector[29])
		data_out <= r_63_29;
		if (write_en==1'b1)
			r_63_29 <= data_in;
	if (addr_selector[63]&addr_selector[30])
		data_out <= r_63_30;
		if (write_en==1'b1)
			r_63_30 <= data_in;
	if (addr_selector[63]&addr_selector[31])
		data_out <= r_63_31;
		if (write_en==1'b1)
			r_63_31 <= data_in;
	if (addr_selector[63]&addr_selector[32])
		data_out <= r_63_32;
		if (write_en==1'b1)
			r_63_32 <= data_in;
	if (addr_selector[63]&addr_selector[33])
		data_out <= r_63_33;
		if (write_en==1'b1)
			r_63_33 <= data_in;
	if (addr_selector[63]&addr_selector[34])
		data_out <= r_63_34;
		if (write_en==1'b1)
			r_63_34 <= data_in;
	if (addr_selector[63]&addr_selector[35])
		data_out <= r_63_35;
		if (write_en==1'b1)
			r_63_35 <= data_in;
	if (addr_selector[63]&addr_selector[36])
		data_out <= r_63_36;
		if (write_en==1'b1)
			r_63_36 <= data_in;
	if (addr_selector[63]&addr_selector[37])
		data_out <= r_63_37;
		if (write_en==1'b1)
			r_63_37 <= data_in;
	if (addr_selector[63]&addr_selector[38])
		data_out <= r_63_38;
		if (write_en==1'b1)
			r_63_38 <= data_in;
	if (addr_selector[63]&addr_selector[39])
		data_out <= r_63_39;
		if (write_en==1'b1)
			r_63_39 <= data_in;
	if (addr_selector[63]&addr_selector[40])
		data_out <= r_63_40;
		if (write_en==1'b1)
			r_63_40 <= data_in;
	if (addr_selector[63]&addr_selector[41])
		data_out <= r_63_41;
		if (write_en==1'b1)
			r_63_41 <= data_in;
	if (addr_selector[63]&addr_selector[42])
		data_out <= r_63_42;
		if (write_en==1'b1)
			r_63_42 <= data_in;
	if (addr_selector[63]&addr_selector[43])
		data_out <= r_63_43;
		if (write_en==1'b1)
			r_63_43 <= data_in;
	if (addr_selector[63]&addr_selector[44])
		data_out <= r_63_44;
		if (write_en==1'b1)
			r_63_44 <= data_in;
	if (addr_selector[63]&addr_selector[45])
		data_out <= r_63_45;
		if (write_en==1'b1)
			r_63_45 <= data_in;
	if (addr_selector[63]&addr_selector[46])
		data_out <= r_63_46;
		if (write_en==1'b1)
			r_63_46 <= data_in;
	if (addr_selector[63]&addr_selector[47])
		data_out <= r_63_47;
		if (write_en==1'b1)
			r_63_47 <= data_in;
	if (addr_selector[63]&addr_selector[48])
		data_out <= r_63_48;
		if (write_en==1'b1)
			r_63_48 <= data_in;
	if (addr_selector[63]&addr_selector[49])
		data_out <= r_63_49;
		if (write_en==1'b1)
			r_63_49 <= data_in;
	if (addr_selector[63]&addr_selector[50])
		data_out <= r_63_50;
		if (write_en==1'b1)
			r_63_50 <= data_in;
	if (addr_selector[63]&addr_selector[51])
		data_out <= r_63_51;
		if (write_en==1'b1)
			r_63_51 <= data_in;
	if (addr_selector[63]&addr_selector[52])
		data_out <= r_63_52;
		if (write_en==1'b1)
			r_63_52 <= data_in;
	if (addr_selector[63]&addr_selector[53])
		data_out <= r_63_53;
		if (write_en==1'b1)
			r_63_53 <= data_in;
	if (addr_selector[63]&addr_selector[54])
		data_out <= r_63_54;
		if (write_en==1'b1)
			r_63_54 <= data_in;
	if (addr_selector[63]&addr_selector[55])
		data_out <= r_63_55;
		if (write_en==1'b1)
			r_63_55 <= data_in;
	if (addr_selector[63]&addr_selector[56])
		data_out <= r_63_56;
		if (write_en==1'b1)
			r_63_56 <= data_in;
	if (addr_selector[63]&addr_selector[57])
		data_out <= r_63_57;
		if (write_en==1'b1)
			r_63_57 <= data_in;
	if (addr_selector[63]&addr_selector[58])
		data_out <= r_63_58;
		if (write_en==1'b1)
			r_63_58 <= data_in;
	if (addr_selector[63]&addr_selector[59])
		data_out <= r_63_59;
		if (write_en==1'b1)
			r_63_59 <= data_in;
	if (addr_selector[63]&addr_selector[60])
		data_out <= r_63_60;
		if (write_en==1'b1)
			r_63_60 <= data_in;
	if (addr_selector[63]&addr_selector[61])
		data_out <= r_63_61;
		if (write_en==1'b1)
			r_63_61 <= data_in;
	if (addr_selector[63]&addr_selector[62])
		data_out <= r_63_62;
		if (write_en==1'b1)
			r_63_62 <= data_in;
	if (addr_selector[63]&addr_selector[63])
		data_out <= r_63_63;
		if (write_en==1'b1)
			r_63_63 <= data_in;
end

endmodule
