module address_decode_12_4
(
input wire[11:0] addr_raw,
output wire[4095:0] addr_selector
);

wire[16:0] r_0_addr;
wire[16:0] r_1_addr;
wire[16:0] r_2_addr;

assign r_0_addr[0] = (addr_raw[3:0]==4'b0000) ?1'b1:1'b0;
assign r_0_addr[1] = (addr_raw[3:0]==4'b0001) ?1'b1:1'b0;
assign r_0_addr[2] = (addr_raw[3:0]==4'b0010) ?1'b1:1'b0;
assign r_0_addr[3] = (addr_raw[3:0]==4'b0011) ?1'b1:1'b0;
assign r_0_addr[4] = (addr_raw[3:0]==4'b0100) ?1'b1:1'b0;
assign r_0_addr[5] = (addr_raw[3:0]==4'b0101) ?1'b1:1'b0;
assign r_0_addr[6] = (addr_raw[3:0]==4'b0110) ?1'b1:1'b0;
assign r_0_addr[7] = (addr_raw[3:0]==4'b0111) ?1'b1:1'b0;
assign r_0_addr[8] = (addr_raw[3:0]==4'b1000) ?1'b1:1'b0;
assign r_0_addr[9] = (addr_raw[3:0]==4'b1001) ?1'b1:1'b0;
assign r_0_addr[10] = (addr_raw[3:0]==4'b1010) ?1'b1:1'b0;
assign r_0_addr[11] = (addr_raw[3:0]==4'b1011) ?1'b1:1'b0;
assign r_0_addr[12] = (addr_raw[3:0]==4'b1100) ?1'b1:1'b0;
assign r_0_addr[13] = (addr_raw[3:0]==4'b1101) ?1'b1:1'b0;
assign r_0_addr[14] = (addr_raw[3:0]==4'b1110) ?1'b1:1'b0;
assign r_0_addr[15] = (addr_raw[3:0]==4'b1111) ?1'b1:1'b0;
assign r_1_addr[0] = (addr_raw[7:4]==4'b0000) ?1'b1:1'b0;
assign r_1_addr[1] = (addr_raw[7:4]==4'b0001) ?1'b1:1'b0;
assign r_1_addr[2] = (addr_raw[7:4]==4'b0010) ?1'b1:1'b0;
assign r_1_addr[3] = (addr_raw[7:4]==4'b0011) ?1'b1:1'b0;
assign r_1_addr[4] = (addr_raw[7:4]==4'b0100) ?1'b1:1'b0;
assign r_1_addr[5] = (addr_raw[7:4]==4'b0101) ?1'b1:1'b0;
assign r_1_addr[6] = (addr_raw[7:4]==4'b0110) ?1'b1:1'b0;
assign r_1_addr[7] = (addr_raw[7:4]==4'b0111) ?1'b1:1'b0;
assign r_1_addr[8] = (addr_raw[7:4]==4'b1000) ?1'b1:1'b0;
assign r_1_addr[9] = (addr_raw[7:4]==4'b1001) ?1'b1:1'b0;
assign r_1_addr[10] = (addr_raw[7:4]==4'b1010) ?1'b1:1'b0;
assign r_1_addr[11] = (addr_raw[7:4]==4'b1011) ?1'b1:1'b0;
assign r_1_addr[12] = (addr_raw[7:4]==4'b1100) ?1'b1:1'b0;
assign r_1_addr[13] = (addr_raw[7:4]==4'b1101) ?1'b1:1'b0;
assign r_1_addr[14] = (addr_raw[7:4]==4'b1110) ?1'b1:1'b0;
assign r_1_addr[15] = (addr_raw[7:4]==4'b1111) ?1'b1:1'b0;
assign r_2_addr[0] = (addr_raw[11:8]==4'b0000) ?1'b1:1'b0;
assign r_2_addr[1] = (addr_raw[11:8]==4'b0001) ?1'b1:1'b0;
assign r_2_addr[2] = (addr_raw[11:8]==4'b0010) ?1'b1:1'b0;
assign r_2_addr[3] = (addr_raw[11:8]==4'b0011) ?1'b1:1'b0;
assign r_2_addr[4] = (addr_raw[11:8]==4'b0100) ?1'b1:1'b0;
assign r_2_addr[5] = (addr_raw[11:8]==4'b0101) ?1'b1:1'b0;
assign r_2_addr[6] = (addr_raw[11:8]==4'b0110) ?1'b1:1'b0;
assign r_2_addr[7] = (addr_raw[11:8]==4'b0111) ?1'b1:1'b0;
assign r_2_addr[8] = (addr_raw[11:8]==4'b1000) ?1'b1:1'b0;
assign r_2_addr[9] = (addr_raw[11:8]==4'b1001) ?1'b1:1'b0;
assign r_2_addr[10] = (addr_raw[11:8]==4'b1010) ?1'b1:1'b0;
assign r_2_addr[11] = (addr_raw[11:8]==4'b1011) ?1'b1:1'b0;
assign r_2_addr[12] = (addr_raw[11:8]==4'b1100) ?1'b1:1'b0;
assign r_2_addr[13] = (addr_raw[11:8]==4'b1101) ?1'b1:1'b0;
assign r_2_addr[14] = (addr_raw[11:8]==4'b1110) ?1'b1:1'b0;
assign r_2_addr[15] = (addr_raw[11:8]==4'b1111) ?1'b1:1'b0;

addr_selector = {r_2_addr[15]&r_1_addr[15]&r_0_addr[15],
r_2_addr[15]&r_1_addr[15]&r_0_addr[14],
r_2_addr[15]&r_1_addr[15]&r_0_addr[13],
r_2_addr[15]&r_1_addr[15]&r_0_addr[12],
r_2_addr[15]&r_1_addr[15]&r_0_addr[11],
r_2_addr[15]&r_1_addr[15]&r_0_addr[10],
r_2_addr[15]&r_1_addr[15]&r_0_addr[9],
r_2_addr[15]&r_1_addr[15]&r_0_addr[8],
r_2_addr[15]&r_1_addr[15]&r_0_addr[7],
r_2_addr[15]&r_1_addr[15]&r_0_addr[6],
r_2_addr[15]&r_1_addr[15]&r_0_addr[5],
r_2_addr[15]&r_1_addr[15]&r_0_addr[4],
r_2_addr[15]&r_1_addr[15]&r_0_addr[3],
r_2_addr[15]&r_1_addr[15]&r_0_addr[2],
r_2_addr[15]&r_1_addr[15]&r_0_addr[1],
r_2_addr[15]&r_1_addr[15]&r_0_addr[0],
r_2_addr[15]&r_1_addr[14]&r_0_addr[15],
r_2_addr[15]&r_1_addr[14]&r_0_addr[14],
r_2_addr[15]&r_1_addr[14]&r_0_addr[13],
r_2_addr[15]&r_1_addr[14]&r_0_addr[12],
r_2_addr[15]&r_1_addr[14]&r_0_addr[11],
r_2_addr[15]&r_1_addr[14]&r_0_addr[10],
r_2_addr[15]&r_1_addr[14]&r_0_addr[9],
r_2_addr[15]&r_1_addr[14]&r_0_addr[8],
r_2_addr[15]&r_1_addr[14]&r_0_addr[7],
r_2_addr[15]&r_1_addr[14]&r_0_addr[6],
r_2_addr[15]&r_1_addr[14]&r_0_addr[5],
r_2_addr[15]&r_1_addr[14]&r_0_addr[4],
r_2_addr[15]&r_1_addr[14]&r_0_addr[3],
r_2_addr[15]&r_1_addr[14]&r_0_addr[2],
r_2_addr[15]&r_1_addr[14]&r_0_addr[1],
r_2_addr[15]&r_1_addr[14]&r_0_addr[0],
r_2_addr[15]&r_1_addr[13]&r_0_addr[15],
r_2_addr[15]&r_1_addr[13]&r_0_addr[14],
r_2_addr[15]&r_1_addr[13]&r_0_addr[13],
r_2_addr[15]&r_1_addr[13]&r_0_addr[12],
r_2_addr[15]&r_1_addr[13]&r_0_addr[11],
r_2_addr[15]&r_1_addr[13]&r_0_addr[10],
r_2_addr[15]&r_1_addr[13]&r_0_addr[9],
r_2_addr[15]&r_1_addr[13]&r_0_addr[8],
r_2_addr[15]&r_1_addr[13]&r_0_addr[7],
r_2_addr[15]&r_1_addr[13]&r_0_addr[6],
r_2_addr[15]&r_1_addr[13]&r_0_addr[5],
r_2_addr[15]&r_1_addr[13]&r_0_addr[4],
r_2_addr[15]&r_1_addr[13]&r_0_addr[3],
r_2_addr[15]&r_1_addr[13]&r_0_addr[2],
r_2_addr[15]&r_1_addr[13]&r_0_addr[1],
r_2_addr[15]&r_1_addr[13]&r_0_addr[0],
r_2_addr[15]&r_1_addr[12]&r_0_addr[15],
r_2_addr[15]&r_1_addr[12]&r_0_addr[14],
r_2_addr[15]&r_1_addr[12]&r_0_addr[13],
r_2_addr[15]&r_1_addr[12]&r_0_addr[12],
r_2_addr[15]&r_1_addr[12]&r_0_addr[11],
r_2_addr[15]&r_1_addr[12]&r_0_addr[10],
r_2_addr[15]&r_1_addr[12]&r_0_addr[9],
r_2_addr[15]&r_1_addr[12]&r_0_addr[8],
r_2_addr[15]&r_1_addr[12]&r_0_addr[7],
r_2_addr[15]&r_1_addr[12]&r_0_addr[6],
r_2_addr[15]&r_1_addr[12]&r_0_addr[5],
r_2_addr[15]&r_1_addr[12]&r_0_addr[4],
r_2_addr[15]&r_1_addr[12]&r_0_addr[3],
r_2_addr[15]&r_1_addr[12]&r_0_addr[2],
r_2_addr[15]&r_1_addr[12]&r_0_addr[1],
r_2_addr[15]&r_1_addr[12]&r_0_addr[0],
r_2_addr[15]&r_1_addr[11]&r_0_addr[15],
r_2_addr[15]&r_1_addr[11]&r_0_addr[14],
r_2_addr[15]&r_1_addr[11]&r_0_addr[13],
r_2_addr[15]&r_1_addr[11]&r_0_addr[12],
r_2_addr[15]&r_1_addr[11]&r_0_addr[11],
r_2_addr[15]&r_1_addr[11]&r_0_addr[10],
r_2_addr[15]&r_1_addr[11]&r_0_addr[9],
r_2_addr[15]&r_1_addr[11]&r_0_addr[8],
r_2_addr[15]&r_1_addr[11]&r_0_addr[7],
r_2_addr[15]&r_1_addr[11]&r_0_addr[6],
r_2_addr[15]&r_1_addr[11]&r_0_addr[5],
r_2_addr[15]&r_1_addr[11]&r_0_addr[4],
r_2_addr[15]&r_1_addr[11]&r_0_addr[3],
r_2_addr[15]&r_1_addr[11]&r_0_addr[2],
r_2_addr[15]&r_1_addr[11]&r_0_addr[1],
r_2_addr[15]&r_1_addr[11]&r_0_addr[0],
r_2_addr[15]&r_1_addr[10]&r_0_addr[15],
r_2_addr[15]&r_1_addr[10]&r_0_addr[14],
r_2_addr[15]&r_1_addr[10]&r_0_addr[13],
r_2_addr[15]&r_1_addr[10]&r_0_addr[12],
r_2_addr[15]&r_1_addr[10]&r_0_addr[11],
r_2_addr[15]&r_1_addr[10]&r_0_addr[10],
r_2_addr[15]&r_1_addr[10]&r_0_addr[9],
r_2_addr[15]&r_1_addr[10]&r_0_addr[8],
r_2_addr[15]&r_1_addr[10]&r_0_addr[7],
r_2_addr[15]&r_1_addr[10]&r_0_addr[6],
r_2_addr[15]&r_1_addr[10]&r_0_addr[5],
r_2_addr[15]&r_1_addr[10]&r_0_addr[4],
r_2_addr[15]&r_1_addr[10]&r_0_addr[3],
r_2_addr[15]&r_1_addr[10]&r_0_addr[2],
r_2_addr[15]&r_1_addr[10]&r_0_addr[1],
r_2_addr[15]&r_1_addr[10]&r_0_addr[0],
r_2_addr[15]&r_1_addr[9]&r_0_addr[15],
r_2_addr[15]&r_1_addr[9]&r_0_addr[14],
r_2_addr[15]&r_1_addr[9]&r_0_addr[13],
r_2_addr[15]&r_1_addr[9]&r_0_addr[12],
r_2_addr[15]&r_1_addr[9]&r_0_addr[11],
r_2_addr[15]&r_1_addr[9]&r_0_addr[10],
r_2_addr[15]&r_1_addr[9]&r_0_addr[9],
r_2_addr[15]&r_1_addr[9]&r_0_addr[8],
r_2_addr[15]&r_1_addr[9]&r_0_addr[7],
r_2_addr[15]&r_1_addr[9]&r_0_addr[6],
r_2_addr[15]&r_1_addr[9]&r_0_addr[5],
r_2_addr[15]&r_1_addr[9]&r_0_addr[4],
r_2_addr[15]&r_1_addr[9]&r_0_addr[3],
r_2_addr[15]&r_1_addr[9]&r_0_addr[2],
r_2_addr[15]&r_1_addr[9]&r_0_addr[1],
r_2_addr[15]&r_1_addr[9]&r_0_addr[0],
r_2_addr[15]&r_1_addr[8]&r_0_addr[15],
r_2_addr[15]&r_1_addr[8]&r_0_addr[14],
r_2_addr[15]&r_1_addr[8]&r_0_addr[13],
r_2_addr[15]&r_1_addr[8]&r_0_addr[12],
r_2_addr[15]&r_1_addr[8]&r_0_addr[11],
r_2_addr[15]&r_1_addr[8]&r_0_addr[10],
r_2_addr[15]&r_1_addr[8]&r_0_addr[9],
r_2_addr[15]&r_1_addr[8]&r_0_addr[8],
r_2_addr[15]&r_1_addr[8]&r_0_addr[7],
r_2_addr[15]&r_1_addr[8]&r_0_addr[6],
r_2_addr[15]&r_1_addr[8]&r_0_addr[5],
r_2_addr[15]&r_1_addr[8]&r_0_addr[4],
r_2_addr[15]&r_1_addr[8]&r_0_addr[3],
r_2_addr[15]&r_1_addr[8]&r_0_addr[2],
r_2_addr[15]&r_1_addr[8]&r_0_addr[1],
r_2_addr[15]&r_1_addr[8]&r_0_addr[0],
r_2_addr[15]&r_1_addr[7]&r_0_addr[15],
r_2_addr[15]&r_1_addr[7]&r_0_addr[14],
r_2_addr[15]&r_1_addr[7]&r_0_addr[13],
r_2_addr[15]&r_1_addr[7]&r_0_addr[12],
r_2_addr[15]&r_1_addr[7]&r_0_addr[11],
r_2_addr[15]&r_1_addr[7]&r_0_addr[10],
r_2_addr[15]&r_1_addr[7]&r_0_addr[9],
r_2_addr[15]&r_1_addr[7]&r_0_addr[8],
r_2_addr[15]&r_1_addr[7]&r_0_addr[7],
r_2_addr[15]&r_1_addr[7]&r_0_addr[6],
r_2_addr[15]&r_1_addr[7]&r_0_addr[5],
r_2_addr[15]&r_1_addr[7]&r_0_addr[4],
r_2_addr[15]&r_1_addr[7]&r_0_addr[3],
r_2_addr[15]&r_1_addr[7]&r_0_addr[2],
r_2_addr[15]&r_1_addr[7]&r_0_addr[1],
r_2_addr[15]&r_1_addr[7]&r_0_addr[0],
r_2_addr[15]&r_1_addr[6]&r_0_addr[15],
r_2_addr[15]&r_1_addr[6]&r_0_addr[14],
r_2_addr[15]&r_1_addr[6]&r_0_addr[13],
r_2_addr[15]&r_1_addr[6]&r_0_addr[12],
r_2_addr[15]&r_1_addr[6]&r_0_addr[11],
r_2_addr[15]&r_1_addr[6]&r_0_addr[10],
r_2_addr[15]&r_1_addr[6]&r_0_addr[9],
r_2_addr[15]&r_1_addr[6]&r_0_addr[8],
r_2_addr[15]&r_1_addr[6]&r_0_addr[7],
r_2_addr[15]&r_1_addr[6]&r_0_addr[6],
r_2_addr[15]&r_1_addr[6]&r_0_addr[5],
r_2_addr[15]&r_1_addr[6]&r_0_addr[4],
r_2_addr[15]&r_1_addr[6]&r_0_addr[3],
r_2_addr[15]&r_1_addr[6]&r_0_addr[2],
r_2_addr[15]&r_1_addr[6]&r_0_addr[1],
r_2_addr[15]&r_1_addr[6]&r_0_addr[0],
r_2_addr[15]&r_1_addr[5]&r_0_addr[15],
r_2_addr[15]&r_1_addr[5]&r_0_addr[14],
r_2_addr[15]&r_1_addr[5]&r_0_addr[13],
r_2_addr[15]&r_1_addr[5]&r_0_addr[12],
r_2_addr[15]&r_1_addr[5]&r_0_addr[11],
r_2_addr[15]&r_1_addr[5]&r_0_addr[10],
r_2_addr[15]&r_1_addr[5]&r_0_addr[9],
r_2_addr[15]&r_1_addr[5]&r_0_addr[8],
r_2_addr[15]&r_1_addr[5]&r_0_addr[7],
r_2_addr[15]&r_1_addr[5]&r_0_addr[6],
r_2_addr[15]&r_1_addr[5]&r_0_addr[5],
r_2_addr[15]&r_1_addr[5]&r_0_addr[4],
r_2_addr[15]&r_1_addr[5]&r_0_addr[3],
r_2_addr[15]&r_1_addr[5]&r_0_addr[2],
r_2_addr[15]&r_1_addr[5]&r_0_addr[1],
r_2_addr[15]&r_1_addr[5]&r_0_addr[0],
r_2_addr[15]&r_1_addr[4]&r_0_addr[15],
r_2_addr[15]&r_1_addr[4]&r_0_addr[14],
r_2_addr[15]&r_1_addr[4]&r_0_addr[13],
r_2_addr[15]&r_1_addr[4]&r_0_addr[12],
r_2_addr[15]&r_1_addr[4]&r_0_addr[11],
r_2_addr[15]&r_1_addr[4]&r_0_addr[10],
r_2_addr[15]&r_1_addr[4]&r_0_addr[9],
r_2_addr[15]&r_1_addr[4]&r_0_addr[8],
r_2_addr[15]&r_1_addr[4]&r_0_addr[7],
r_2_addr[15]&r_1_addr[4]&r_0_addr[6],
r_2_addr[15]&r_1_addr[4]&r_0_addr[5],
r_2_addr[15]&r_1_addr[4]&r_0_addr[4],
r_2_addr[15]&r_1_addr[4]&r_0_addr[3],
r_2_addr[15]&r_1_addr[4]&r_0_addr[2],
r_2_addr[15]&r_1_addr[4]&r_0_addr[1],
r_2_addr[15]&r_1_addr[4]&r_0_addr[0],
r_2_addr[15]&r_1_addr[3]&r_0_addr[15],
r_2_addr[15]&r_1_addr[3]&r_0_addr[14],
r_2_addr[15]&r_1_addr[3]&r_0_addr[13],
r_2_addr[15]&r_1_addr[3]&r_0_addr[12],
r_2_addr[15]&r_1_addr[3]&r_0_addr[11],
r_2_addr[15]&r_1_addr[3]&r_0_addr[10],
r_2_addr[15]&r_1_addr[3]&r_0_addr[9],
r_2_addr[15]&r_1_addr[3]&r_0_addr[8],
r_2_addr[15]&r_1_addr[3]&r_0_addr[7],
r_2_addr[15]&r_1_addr[3]&r_0_addr[6],
r_2_addr[15]&r_1_addr[3]&r_0_addr[5],
r_2_addr[15]&r_1_addr[3]&r_0_addr[4],
r_2_addr[15]&r_1_addr[3]&r_0_addr[3],
r_2_addr[15]&r_1_addr[3]&r_0_addr[2],
r_2_addr[15]&r_1_addr[3]&r_0_addr[1],
r_2_addr[15]&r_1_addr[3]&r_0_addr[0],
r_2_addr[15]&r_1_addr[2]&r_0_addr[15],
r_2_addr[15]&r_1_addr[2]&r_0_addr[14],
r_2_addr[15]&r_1_addr[2]&r_0_addr[13],
r_2_addr[15]&r_1_addr[2]&r_0_addr[12],
r_2_addr[15]&r_1_addr[2]&r_0_addr[11],
r_2_addr[15]&r_1_addr[2]&r_0_addr[10],
r_2_addr[15]&r_1_addr[2]&r_0_addr[9],
r_2_addr[15]&r_1_addr[2]&r_0_addr[8],
r_2_addr[15]&r_1_addr[2]&r_0_addr[7],
r_2_addr[15]&r_1_addr[2]&r_0_addr[6],
r_2_addr[15]&r_1_addr[2]&r_0_addr[5],
r_2_addr[15]&r_1_addr[2]&r_0_addr[4],
r_2_addr[15]&r_1_addr[2]&r_0_addr[3],
r_2_addr[15]&r_1_addr[2]&r_0_addr[2],
r_2_addr[15]&r_1_addr[2]&r_0_addr[1],
r_2_addr[15]&r_1_addr[2]&r_0_addr[0],
r_2_addr[15]&r_1_addr[1]&r_0_addr[15],
r_2_addr[15]&r_1_addr[1]&r_0_addr[14],
r_2_addr[15]&r_1_addr[1]&r_0_addr[13],
r_2_addr[15]&r_1_addr[1]&r_0_addr[12],
r_2_addr[15]&r_1_addr[1]&r_0_addr[11],
r_2_addr[15]&r_1_addr[1]&r_0_addr[10],
r_2_addr[15]&r_1_addr[1]&r_0_addr[9],
r_2_addr[15]&r_1_addr[1]&r_0_addr[8],
r_2_addr[15]&r_1_addr[1]&r_0_addr[7],
r_2_addr[15]&r_1_addr[1]&r_0_addr[6],
r_2_addr[15]&r_1_addr[1]&r_0_addr[5],
r_2_addr[15]&r_1_addr[1]&r_0_addr[4],
r_2_addr[15]&r_1_addr[1]&r_0_addr[3],
r_2_addr[15]&r_1_addr[1]&r_0_addr[2],
r_2_addr[15]&r_1_addr[1]&r_0_addr[1],
r_2_addr[15]&r_1_addr[1]&r_0_addr[0],
r_2_addr[15]&r_1_addr[0]&r_0_addr[15],
r_2_addr[15]&r_1_addr[0]&r_0_addr[14],
r_2_addr[15]&r_1_addr[0]&r_0_addr[13],
r_2_addr[15]&r_1_addr[0]&r_0_addr[12],
r_2_addr[15]&r_1_addr[0]&r_0_addr[11],
r_2_addr[15]&r_1_addr[0]&r_0_addr[10],
r_2_addr[15]&r_1_addr[0]&r_0_addr[9],
r_2_addr[15]&r_1_addr[0]&r_0_addr[8],
r_2_addr[15]&r_1_addr[0]&r_0_addr[7],
r_2_addr[15]&r_1_addr[0]&r_0_addr[6],
r_2_addr[15]&r_1_addr[0]&r_0_addr[5],
r_2_addr[15]&r_1_addr[0]&r_0_addr[4],
r_2_addr[15]&r_1_addr[0]&r_0_addr[3],
r_2_addr[15]&r_1_addr[0]&r_0_addr[2],
r_2_addr[15]&r_1_addr[0]&r_0_addr[1],
r_2_addr[15]&r_1_addr[0]&r_0_addr[0],
r_2_addr[14]&r_1_addr[15]&r_0_addr[15],
r_2_addr[14]&r_1_addr[15]&r_0_addr[14],
r_2_addr[14]&r_1_addr[15]&r_0_addr[13],
r_2_addr[14]&r_1_addr[15]&r_0_addr[12],
r_2_addr[14]&r_1_addr[15]&r_0_addr[11],
r_2_addr[14]&r_1_addr[15]&r_0_addr[10],
r_2_addr[14]&r_1_addr[15]&r_0_addr[9],
r_2_addr[14]&r_1_addr[15]&r_0_addr[8],
r_2_addr[14]&r_1_addr[15]&r_0_addr[7],
r_2_addr[14]&r_1_addr[15]&r_0_addr[6],
r_2_addr[14]&r_1_addr[15]&r_0_addr[5],
r_2_addr[14]&r_1_addr[15]&r_0_addr[4],
r_2_addr[14]&r_1_addr[15]&r_0_addr[3],
r_2_addr[14]&r_1_addr[15]&r_0_addr[2],
r_2_addr[14]&r_1_addr[15]&r_0_addr[1],
r_2_addr[14]&r_1_addr[15]&r_0_addr[0],
r_2_addr[14]&r_1_addr[14]&r_0_addr[15],
r_2_addr[14]&r_1_addr[14]&r_0_addr[14],
r_2_addr[14]&r_1_addr[14]&r_0_addr[13],
r_2_addr[14]&r_1_addr[14]&r_0_addr[12],
r_2_addr[14]&r_1_addr[14]&r_0_addr[11],
r_2_addr[14]&r_1_addr[14]&r_0_addr[10],
r_2_addr[14]&r_1_addr[14]&r_0_addr[9],
r_2_addr[14]&r_1_addr[14]&r_0_addr[8],
r_2_addr[14]&r_1_addr[14]&r_0_addr[7],
r_2_addr[14]&r_1_addr[14]&r_0_addr[6],
r_2_addr[14]&r_1_addr[14]&r_0_addr[5],
r_2_addr[14]&r_1_addr[14]&r_0_addr[4],
r_2_addr[14]&r_1_addr[14]&r_0_addr[3],
r_2_addr[14]&r_1_addr[14]&r_0_addr[2],
r_2_addr[14]&r_1_addr[14]&r_0_addr[1],
r_2_addr[14]&r_1_addr[14]&r_0_addr[0],
r_2_addr[14]&r_1_addr[13]&r_0_addr[15],
r_2_addr[14]&r_1_addr[13]&r_0_addr[14],
r_2_addr[14]&r_1_addr[13]&r_0_addr[13],
r_2_addr[14]&r_1_addr[13]&r_0_addr[12],
r_2_addr[14]&r_1_addr[13]&r_0_addr[11],
r_2_addr[14]&r_1_addr[13]&r_0_addr[10],
r_2_addr[14]&r_1_addr[13]&r_0_addr[9],
r_2_addr[14]&r_1_addr[13]&r_0_addr[8],
r_2_addr[14]&r_1_addr[13]&r_0_addr[7],
r_2_addr[14]&r_1_addr[13]&r_0_addr[6],
r_2_addr[14]&r_1_addr[13]&r_0_addr[5],
r_2_addr[14]&r_1_addr[13]&r_0_addr[4],
r_2_addr[14]&r_1_addr[13]&r_0_addr[3],
r_2_addr[14]&r_1_addr[13]&r_0_addr[2],
r_2_addr[14]&r_1_addr[13]&r_0_addr[1],
r_2_addr[14]&r_1_addr[13]&r_0_addr[0],
r_2_addr[14]&r_1_addr[12]&r_0_addr[15],
r_2_addr[14]&r_1_addr[12]&r_0_addr[14],
r_2_addr[14]&r_1_addr[12]&r_0_addr[13],
r_2_addr[14]&r_1_addr[12]&r_0_addr[12],
r_2_addr[14]&r_1_addr[12]&r_0_addr[11],
r_2_addr[14]&r_1_addr[12]&r_0_addr[10],
r_2_addr[14]&r_1_addr[12]&r_0_addr[9],
r_2_addr[14]&r_1_addr[12]&r_0_addr[8],
r_2_addr[14]&r_1_addr[12]&r_0_addr[7],
r_2_addr[14]&r_1_addr[12]&r_0_addr[6],
r_2_addr[14]&r_1_addr[12]&r_0_addr[5],
r_2_addr[14]&r_1_addr[12]&r_0_addr[4],
r_2_addr[14]&r_1_addr[12]&r_0_addr[3],
r_2_addr[14]&r_1_addr[12]&r_0_addr[2],
r_2_addr[14]&r_1_addr[12]&r_0_addr[1],
r_2_addr[14]&r_1_addr[12]&r_0_addr[0],
r_2_addr[14]&r_1_addr[11]&r_0_addr[15],
r_2_addr[14]&r_1_addr[11]&r_0_addr[14],
r_2_addr[14]&r_1_addr[11]&r_0_addr[13],
r_2_addr[14]&r_1_addr[11]&r_0_addr[12],
r_2_addr[14]&r_1_addr[11]&r_0_addr[11],
r_2_addr[14]&r_1_addr[11]&r_0_addr[10],
r_2_addr[14]&r_1_addr[11]&r_0_addr[9],
r_2_addr[14]&r_1_addr[11]&r_0_addr[8],
r_2_addr[14]&r_1_addr[11]&r_0_addr[7],
r_2_addr[14]&r_1_addr[11]&r_0_addr[6],
r_2_addr[14]&r_1_addr[11]&r_0_addr[5],
r_2_addr[14]&r_1_addr[11]&r_0_addr[4],
r_2_addr[14]&r_1_addr[11]&r_0_addr[3],
r_2_addr[14]&r_1_addr[11]&r_0_addr[2],
r_2_addr[14]&r_1_addr[11]&r_0_addr[1],
r_2_addr[14]&r_1_addr[11]&r_0_addr[0],
r_2_addr[14]&r_1_addr[10]&r_0_addr[15],
r_2_addr[14]&r_1_addr[10]&r_0_addr[14],
r_2_addr[14]&r_1_addr[10]&r_0_addr[13],
r_2_addr[14]&r_1_addr[10]&r_0_addr[12],
r_2_addr[14]&r_1_addr[10]&r_0_addr[11],
r_2_addr[14]&r_1_addr[10]&r_0_addr[10],
r_2_addr[14]&r_1_addr[10]&r_0_addr[9],
r_2_addr[14]&r_1_addr[10]&r_0_addr[8],
r_2_addr[14]&r_1_addr[10]&r_0_addr[7],
r_2_addr[14]&r_1_addr[10]&r_0_addr[6],
r_2_addr[14]&r_1_addr[10]&r_0_addr[5],
r_2_addr[14]&r_1_addr[10]&r_0_addr[4],
r_2_addr[14]&r_1_addr[10]&r_0_addr[3],
r_2_addr[14]&r_1_addr[10]&r_0_addr[2],
r_2_addr[14]&r_1_addr[10]&r_0_addr[1],
r_2_addr[14]&r_1_addr[10]&r_0_addr[0],
r_2_addr[14]&r_1_addr[9]&r_0_addr[15],
r_2_addr[14]&r_1_addr[9]&r_0_addr[14],
r_2_addr[14]&r_1_addr[9]&r_0_addr[13],
r_2_addr[14]&r_1_addr[9]&r_0_addr[12],
r_2_addr[14]&r_1_addr[9]&r_0_addr[11],
r_2_addr[14]&r_1_addr[9]&r_0_addr[10],
r_2_addr[14]&r_1_addr[9]&r_0_addr[9],
r_2_addr[14]&r_1_addr[9]&r_0_addr[8],
r_2_addr[14]&r_1_addr[9]&r_0_addr[7],
r_2_addr[14]&r_1_addr[9]&r_0_addr[6],
r_2_addr[14]&r_1_addr[9]&r_0_addr[5],
r_2_addr[14]&r_1_addr[9]&r_0_addr[4],
r_2_addr[14]&r_1_addr[9]&r_0_addr[3],
r_2_addr[14]&r_1_addr[9]&r_0_addr[2],
r_2_addr[14]&r_1_addr[9]&r_0_addr[1],
r_2_addr[14]&r_1_addr[9]&r_0_addr[0],
r_2_addr[14]&r_1_addr[8]&r_0_addr[15],
r_2_addr[14]&r_1_addr[8]&r_0_addr[14],
r_2_addr[14]&r_1_addr[8]&r_0_addr[13],
r_2_addr[14]&r_1_addr[8]&r_0_addr[12],
r_2_addr[14]&r_1_addr[8]&r_0_addr[11],
r_2_addr[14]&r_1_addr[8]&r_0_addr[10],
r_2_addr[14]&r_1_addr[8]&r_0_addr[9],
r_2_addr[14]&r_1_addr[8]&r_0_addr[8],
r_2_addr[14]&r_1_addr[8]&r_0_addr[7],
r_2_addr[14]&r_1_addr[8]&r_0_addr[6],
r_2_addr[14]&r_1_addr[8]&r_0_addr[5],
r_2_addr[14]&r_1_addr[8]&r_0_addr[4],
r_2_addr[14]&r_1_addr[8]&r_0_addr[3],
r_2_addr[14]&r_1_addr[8]&r_0_addr[2],
r_2_addr[14]&r_1_addr[8]&r_0_addr[1],
r_2_addr[14]&r_1_addr[8]&r_0_addr[0],
r_2_addr[14]&r_1_addr[7]&r_0_addr[15],
r_2_addr[14]&r_1_addr[7]&r_0_addr[14],
r_2_addr[14]&r_1_addr[7]&r_0_addr[13],
r_2_addr[14]&r_1_addr[7]&r_0_addr[12],
r_2_addr[14]&r_1_addr[7]&r_0_addr[11],
r_2_addr[14]&r_1_addr[7]&r_0_addr[10],
r_2_addr[14]&r_1_addr[7]&r_0_addr[9],
r_2_addr[14]&r_1_addr[7]&r_0_addr[8],
r_2_addr[14]&r_1_addr[7]&r_0_addr[7],
r_2_addr[14]&r_1_addr[7]&r_0_addr[6],
r_2_addr[14]&r_1_addr[7]&r_0_addr[5],
r_2_addr[14]&r_1_addr[7]&r_0_addr[4],
r_2_addr[14]&r_1_addr[7]&r_0_addr[3],
r_2_addr[14]&r_1_addr[7]&r_0_addr[2],
r_2_addr[14]&r_1_addr[7]&r_0_addr[1],
r_2_addr[14]&r_1_addr[7]&r_0_addr[0],
r_2_addr[14]&r_1_addr[6]&r_0_addr[15],
r_2_addr[14]&r_1_addr[6]&r_0_addr[14],
r_2_addr[14]&r_1_addr[6]&r_0_addr[13],
r_2_addr[14]&r_1_addr[6]&r_0_addr[12],
r_2_addr[14]&r_1_addr[6]&r_0_addr[11],
r_2_addr[14]&r_1_addr[6]&r_0_addr[10],
r_2_addr[14]&r_1_addr[6]&r_0_addr[9],
r_2_addr[14]&r_1_addr[6]&r_0_addr[8],
r_2_addr[14]&r_1_addr[6]&r_0_addr[7],
r_2_addr[14]&r_1_addr[6]&r_0_addr[6],
r_2_addr[14]&r_1_addr[6]&r_0_addr[5],
r_2_addr[14]&r_1_addr[6]&r_0_addr[4],
r_2_addr[14]&r_1_addr[6]&r_0_addr[3],
r_2_addr[14]&r_1_addr[6]&r_0_addr[2],
r_2_addr[14]&r_1_addr[6]&r_0_addr[1],
r_2_addr[14]&r_1_addr[6]&r_0_addr[0],
r_2_addr[14]&r_1_addr[5]&r_0_addr[15],
r_2_addr[14]&r_1_addr[5]&r_0_addr[14],
r_2_addr[14]&r_1_addr[5]&r_0_addr[13],
r_2_addr[14]&r_1_addr[5]&r_0_addr[12],
r_2_addr[14]&r_1_addr[5]&r_0_addr[11],
r_2_addr[14]&r_1_addr[5]&r_0_addr[10],
r_2_addr[14]&r_1_addr[5]&r_0_addr[9],
r_2_addr[14]&r_1_addr[5]&r_0_addr[8],
r_2_addr[14]&r_1_addr[5]&r_0_addr[7],
r_2_addr[14]&r_1_addr[5]&r_0_addr[6],
r_2_addr[14]&r_1_addr[5]&r_0_addr[5],
r_2_addr[14]&r_1_addr[5]&r_0_addr[4],
r_2_addr[14]&r_1_addr[5]&r_0_addr[3],
r_2_addr[14]&r_1_addr[5]&r_0_addr[2],
r_2_addr[14]&r_1_addr[5]&r_0_addr[1],
r_2_addr[14]&r_1_addr[5]&r_0_addr[0],
r_2_addr[14]&r_1_addr[4]&r_0_addr[15],
r_2_addr[14]&r_1_addr[4]&r_0_addr[14],
r_2_addr[14]&r_1_addr[4]&r_0_addr[13],
r_2_addr[14]&r_1_addr[4]&r_0_addr[12],
r_2_addr[14]&r_1_addr[4]&r_0_addr[11],
r_2_addr[14]&r_1_addr[4]&r_0_addr[10],
r_2_addr[14]&r_1_addr[4]&r_0_addr[9],
r_2_addr[14]&r_1_addr[4]&r_0_addr[8],
r_2_addr[14]&r_1_addr[4]&r_0_addr[7],
r_2_addr[14]&r_1_addr[4]&r_0_addr[6],
r_2_addr[14]&r_1_addr[4]&r_0_addr[5],
r_2_addr[14]&r_1_addr[4]&r_0_addr[4],
r_2_addr[14]&r_1_addr[4]&r_0_addr[3],
r_2_addr[14]&r_1_addr[4]&r_0_addr[2],
r_2_addr[14]&r_1_addr[4]&r_0_addr[1],
r_2_addr[14]&r_1_addr[4]&r_0_addr[0],
r_2_addr[14]&r_1_addr[3]&r_0_addr[15],
r_2_addr[14]&r_1_addr[3]&r_0_addr[14],
r_2_addr[14]&r_1_addr[3]&r_0_addr[13],
r_2_addr[14]&r_1_addr[3]&r_0_addr[12],
r_2_addr[14]&r_1_addr[3]&r_0_addr[11],
r_2_addr[14]&r_1_addr[3]&r_0_addr[10],
r_2_addr[14]&r_1_addr[3]&r_0_addr[9],
r_2_addr[14]&r_1_addr[3]&r_0_addr[8],
r_2_addr[14]&r_1_addr[3]&r_0_addr[7],
r_2_addr[14]&r_1_addr[3]&r_0_addr[6],
r_2_addr[14]&r_1_addr[3]&r_0_addr[5],
r_2_addr[14]&r_1_addr[3]&r_0_addr[4],
r_2_addr[14]&r_1_addr[3]&r_0_addr[3],
r_2_addr[14]&r_1_addr[3]&r_0_addr[2],
r_2_addr[14]&r_1_addr[3]&r_0_addr[1],
r_2_addr[14]&r_1_addr[3]&r_0_addr[0],
r_2_addr[14]&r_1_addr[2]&r_0_addr[15],
r_2_addr[14]&r_1_addr[2]&r_0_addr[14],
r_2_addr[14]&r_1_addr[2]&r_0_addr[13],
r_2_addr[14]&r_1_addr[2]&r_0_addr[12],
r_2_addr[14]&r_1_addr[2]&r_0_addr[11],
r_2_addr[14]&r_1_addr[2]&r_0_addr[10],
r_2_addr[14]&r_1_addr[2]&r_0_addr[9],
r_2_addr[14]&r_1_addr[2]&r_0_addr[8],
r_2_addr[14]&r_1_addr[2]&r_0_addr[7],
r_2_addr[14]&r_1_addr[2]&r_0_addr[6],
r_2_addr[14]&r_1_addr[2]&r_0_addr[5],
r_2_addr[14]&r_1_addr[2]&r_0_addr[4],
r_2_addr[14]&r_1_addr[2]&r_0_addr[3],
r_2_addr[14]&r_1_addr[2]&r_0_addr[2],
r_2_addr[14]&r_1_addr[2]&r_0_addr[1],
r_2_addr[14]&r_1_addr[2]&r_0_addr[0],
r_2_addr[14]&r_1_addr[1]&r_0_addr[15],
r_2_addr[14]&r_1_addr[1]&r_0_addr[14],
r_2_addr[14]&r_1_addr[1]&r_0_addr[13],
r_2_addr[14]&r_1_addr[1]&r_0_addr[12],
r_2_addr[14]&r_1_addr[1]&r_0_addr[11],
r_2_addr[14]&r_1_addr[1]&r_0_addr[10],
r_2_addr[14]&r_1_addr[1]&r_0_addr[9],
r_2_addr[14]&r_1_addr[1]&r_0_addr[8],
r_2_addr[14]&r_1_addr[1]&r_0_addr[7],
r_2_addr[14]&r_1_addr[1]&r_0_addr[6],
r_2_addr[14]&r_1_addr[1]&r_0_addr[5],
r_2_addr[14]&r_1_addr[1]&r_0_addr[4],
r_2_addr[14]&r_1_addr[1]&r_0_addr[3],
r_2_addr[14]&r_1_addr[1]&r_0_addr[2],
r_2_addr[14]&r_1_addr[1]&r_0_addr[1],
r_2_addr[14]&r_1_addr[1]&r_0_addr[0],
r_2_addr[14]&r_1_addr[0]&r_0_addr[15],
r_2_addr[14]&r_1_addr[0]&r_0_addr[14],
r_2_addr[14]&r_1_addr[0]&r_0_addr[13],
r_2_addr[14]&r_1_addr[0]&r_0_addr[12],
r_2_addr[14]&r_1_addr[0]&r_0_addr[11],
r_2_addr[14]&r_1_addr[0]&r_0_addr[10],
r_2_addr[14]&r_1_addr[0]&r_0_addr[9],
r_2_addr[14]&r_1_addr[0]&r_0_addr[8],
r_2_addr[14]&r_1_addr[0]&r_0_addr[7],
r_2_addr[14]&r_1_addr[0]&r_0_addr[6],
r_2_addr[14]&r_1_addr[0]&r_0_addr[5],
r_2_addr[14]&r_1_addr[0]&r_0_addr[4],
r_2_addr[14]&r_1_addr[0]&r_0_addr[3],
r_2_addr[14]&r_1_addr[0]&r_0_addr[2],
r_2_addr[14]&r_1_addr[0]&r_0_addr[1],
r_2_addr[14]&r_1_addr[0]&r_0_addr[0],
r_2_addr[13]&r_1_addr[15]&r_0_addr[15],
r_2_addr[13]&r_1_addr[15]&r_0_addr[14],
r_2_addr[13]&r_1_addr[15]&r_0_addr[13],
r_2_addr[13]&r_1_addr[15]&r_0_addr[12],
r_2_addr[13]&r_1_addr[15]&r_0_addr[11],
r_2_addr[13]&r_1_addr[15]&r_0_addr[10],
r_2_addr[13]&r_1_addr[15]&r_0_addr[9],
r_2_addr[13]&r_1_addr[15]&r_0_addr[8],
r_2_addr[13]&r_1_addr[15]&r_0_addr[7],
r_2_addr[13]&r_1_addr[15]&r_0_addr[6],
r_2_addr[13]&r_1_addr[15]&r_0_addr[5],
r_2_addr[13]&r_1_addr[15]&r_0_addr[4],
r_2_addr[13]&r_1_addr[15]&r_0_addr[3],
r_2_addr[13]&r_1_addr[15]&r_0_addr[2],
r_2_addr[13]&r_1_addr[15]&r_0_addr[1],
r_2_addr[13]&r_1_addr[15]&r_0_addr[0],
r_2_addr[13]&r_1_addr[14]&r_0_addr[15],
r_2_addr[13]&r_1_addr[14]&r_0_addr[14],
r_2_addr[13]&r_1_addr[14]&r_0_addr[13],
r_2_addr[13]&r_1_addr[14]&r_0_addr[12],
r_2_addr[13]&r_1_addr[14]&r_0_addr[11],
r_2_addr[13]&r_1_addr[14]&r_0_addr[10],
r_2_addr[13]&r_1_addr[14]&r_0_addr[9],
r_2_addr[13]&r_1_addr[14]&r_0_addr[8],
r_2_addr[13]&r_1_addr[14]&r_0_addr[7],
r_2_addr[13]&r_1_addr[14]&r_0_addr[6],
r_2_addr[13]&r_1_addr[14]&r_0_addr[5],
r_2_addr[13]&r_1_addr[14]&r_0_addr[4],
r_2_addr[13]&r_1_addr[14]&r_0_addr[3],
r_2_addr[13]&r_1_addr[14]&r_0_addr[2],
r_2_addr[13]&r_1_addr[14]&r_0_addr[1],
r_2_addr[13]&r_1_addr[14]&r_0_addr[0],
r_2_addr[13]&r_1_addr[13]&r_0_addr[15],
r_2_addr[13]&r_1_addr[13]&r_0_addr[14],
r_2_addr[13]&r_1_addr[13]&r_0_addr[13],
r_2_addr[13]&r_1_addr[13]&r_0_addr[12],
r_2_addr[13]&r_1_addr[13]&r_0_addr[11],
r_2_addr[13]&r_1_addr[13]&r_0_addr[10],
r_2_addr[13]&r_1_addr[13]&r_0_addr[9],
r_2_addr[13]&r_1_addr[13]&r_0_addr[8],
r_2_addr[13]&r_1_addr[13]&r_0_addr[7],
r_2_addr[13]&r_1_addr[13]&r_0_addr[6],
r_2_addr[13]&r_1_addr[13]&r_0_addr[5],
r_2_addr[13]&r_1_addr[13]&r_0_addr[4],
r_2_addr[13]&r_1_addr[13]&r_0_addr[3],
r_2_addr[13]&r_1_addr[13]&r_0_addr[2],
r_2_addr[13]&r_1_addr[13]&r_0_addr[1],
r_2_addr[13]&r_1_addr[13]&r_0_addr[0],
r_2_addr[13]&r_1_addr[12]&r_0_addr[15],
r_2_addr[13]&r_1_addr[12]&r_0_addr[14],
r_2_addr[13]&r_1_addr[12]&r_0_addr[13],
r_2_addr[13]&r_1_addr[12]&r_0_addr[12],
r_2_addr[13]&r_1_addr[12]&r_0_addr[11],
r_2_addr[13]&r_1_addr[12]&r_0_addr[10],
r_2_addr[13]&r_1_addr[12]&r_0_addr[9],
r_2_addr[13]&r_1_addr[12]&r_0_addr[8],
r_2_addr[13]&r_1_addr[12]&r_0_addr[7],
r_2_addr[13]&r_1_addr[12]&r_0_addr[6],
r_2_addr[13]&r_1_addr[12]&r_0_addr[5],
r_2_addr[13]&r_1_addr[12]&r_0_addr[4],
r_2_addr[13]&r_1_addr[12]&r_0_addr[3],
r_2_addr[13]&r_1_addr[12]&r_0_addr[2],
r_2_addr[13]&r_1_addr[12]&r_0_addr[1],
r_2_addr[13]&r_1_addr[12]&r_0_addr[0],
r_2_addr[13]&r_1_addr[11]&r_0_addr[15],
r_2_addr[13]&r_1_addr[11]&r_0_addr[14],
r_2_addr[13]&r_1_addr[11]&r_0_addr[13],
r_2_addr[13]&r_1_addr[11]&r_0_addr[12],
r_2_addr[13]&r_1_addr[11]&r_0_addr[11],
r_2_addr[13]&r_1_addr[11]&r_0_addr[10],
r_2_addr[13]&r_1_addr[11]&r_0_addr[9],
r_2_addr[13]&r_1_addr[11]&r_0_addr[8],
r_2_addr[13]&r_1_addr[11]&r_0_addr[7],
r_2_addr[13]&r_1_addr[11]&r_0_addr[6],
r_2_addr[13]&r_1_addr[11]&r_0_addr[5],
r_2_addr[13]&r_1_addr[11]&r_0_addr[4],
r_2_addr[13]&r_1_addr[11]&r_0_addr[3],
r_2_addr[13]&r_1_addr[11]&r_0_addr[2],
r_2_addr[13]&r_1_addr[11]&r_0_addr[1],
r_2_addr[13]&r_1_addr[11]&r_0_addr[0],
r_2_addr[13]&r_1_addr[10]&r_0_addr[15],
r_2_addr[13]&r_1_addr[10]&r_0_addr[14],
r_2_addr[13]&r_1_addr[10]&r_0_addr[13],
r_2_addr[13]&r_1_addr[10]&r_0_addr[12],
r_2_addr[13]&r_1_addr[10]&r_0_addr[11],
r_2_addr[13]&r_1_addr[10]&r_0_addr[10],
r_2_addr[13]&r_1_addr[10]&r_0_addr[9],
r_2_addr[13]&r_1_addr[10]&r_0_addr[8],
r_2_addr[13]&r_1_addr[10]&r_0_addr[7],
r_2_addr[13]&r_1_addr[10]&r_0_addr[6],
r_2_addr[13]&r_1_addr[10]&r_0_addr[5],
r_2_addr[13]&r_1_addr[10]&r_0_addr[4],
r_2_addr[13]&r_1_addr[10]&r_0_addr[3],
r_2_addr[13]&r_1_addr[10]&r_0_addr[2],
r_2_addr[13]&r_1_addr[10]&r_0_addr[1],
r_2_addr[13]&r_1_addr[10]&r_0_addr[0],
r_2_addr[13]&r_1_addr[9]&r_0_addr[15],
r_2_addr[13]&r_1_addr[9]&r_0_addr[14],
r_2_addr[13]&r_1_addr[9]&r_0_addr[13],
r_2_addr[13]&r_1_addr[9]&r_0_addr[12],
r_2_addr[13]&r_1_addr[9]&r_0_addr[11],
r_2_addr[13]&r_1_addr[9]&r_0_addr[10],
r_2_addr[13]&r_1_addr[9]&r_0_addr[9],
r_2_addr[13]&r_1_addr[9]&r_0_addr[8],
r_2_addr[13]&r_1_addr[9]&r_0_addr[7],
r_2_addr[13]&r_1_addr[9]&r_0_addr[6],
r_2_addr[13]&r_1_addr[9]&r_0_addr[5],
r_2_addr[13]&r_1_addr[9]&r_0_addr[4],
r_2_addr[13]&r_1_addr[9]&r_0_addr[3],
r_2_addr[13]&r_1_addr[9]&r_0_addr[2],
r_2_addr[13]&r_1_addr[9]&r_0_addr[1],
r_2_addr[13]&r_1_addr[9]&r_0_addr[0],
r_2_addr[13]&r_1_addr[8]&r_0_addr[15],
r_2_addr[13]&r_1_addr[8]&r_0_addr[14],
r_2_addr[13]&r_1_addr[8]&r_0_addr[13],
r_2_addr[13]&r_1_addr[8]&r_0_addr[12],
r_2_addr[13]&r_1_addr[8]&r_0_addr[11],
r_2_addr[13]&r_1_addr[8]&r_0_addr[10],
r_2_addr[13]&r_1_addr[8]&r_0_addr[9],
r_2_addr[13]&r_1_addr[8]&r_0_addr[8],
r_2_addr[13]&r_1_addr[8]&r_0_addr[7],
r_2_addr[13]&r_1_addr[8]&r_0_addr[6],
r_2_addr[13]&r_1_addr[8]&r_0_addr[5],
r_2_addr[13]&r_1_addr[8]&r_0_addr[4],
r_2_addr[13]&r_1_addr[8]&r_0_addr[3],
r_2_addr[13]&r_1_addr[8]&r_0_addr[2],
r_2_addr[13]&r_1_addr[8]&r_0_addr[1],
r_2_addr[13]&r_1_addr[8]&r_0_addr[0],
r_2_addr[13]&r_1_addr[7]&r_0_addr[15],
r_2_addr[13]&r_1_addr[7]&r_0_addr[14],
r_2_addr[13]&r_1_addr[7]&r_0_addr[13],
r_2_addr[13]&r_1_addr[7]&r_0_addr[12],
r_2_addr[13]&r_1_addr[7]&r_0_addr[11],
r_2_addr[13]&r_1_addr[7]&r_0_addr[10],
r_2_addr[13]&r_1_addr[7]&r_0_addr[9],
r_2_addr[13]&r_1_addr[7]&r_0_addr[8],
r_2_addr[13]&r_1_addr[7]&r_0_addr[7],
r_2_addr[13]&r_1_addr[7]&r_0_addr[6],
r_2_addr[13]&r_1_addr[7]&r_0_addr[5],
r_2_addr[13]&r_1_addr[7]&r_0_addr[4],
r_2_addr[13]&r_1_addr[7]&r_0_addr[3],
r_2_addr[13]&r_1_addr[7]&r_0_addr[2],
r_2_addr[13]&r_1_addr[7]&r_0_addr[1],
r_2_addr[13]&r_1_addr[7]&r_0_addr[0],
r_2_addr[13]&r_1_addr[6]&r_0_addr[15],
r_2_addr[13]&r_1_addr[6]&r_0_addr[14],
r_2_addr[13]&r_1_addr[6]&r_0_addr[13],
r_2_addr[13]&r_1_addr[6]&r_0_addr[12],
r_2_addr[13]&r_1_addr[6]&r_0_addr[11],
r_2_addr[13]&r_1_addr[6]&r_0_addr[10],
r_2_addr[13]&r_1_addr[6]&r_0_addr[9],
r_2_addr[13]&r_1_addr[6]&r_0_addr[8],
r_2_addr[13]&r_1_addr[6]&r_0_addr[7],
r_2_addr[13]&r_1_addr[6]&r_0_addr[6],
r_2_addr[13]&r_1_addr[6]&r_0_addr[5],
r_2_addr[13]&r_1_addr[6]&r_0_addr[4],
r_2_addr[13]&r_1_addr[6]&r_0_addr[3],
r_2_addr[13]&r_1_addr[6]&r_0_addr[2],
r_2_addr[13]&r_1_addr[6]&r_0_addr[1],
r_2_addr[13]&r_1_addr[6]&r_0_addr[0],
r_2_addr[13]&r_1_addr[5]&r_0_addr[15],
r_2_addr[13]&r_1_addr[5]&r_0_addr[14],
r_2_addr[13]&r_1_addr[5]&r_0_addr[13],
r_2_addr[13]&r_1_addr[5]&r_0_addr[12],
r_2_addr[13]&r_1_addr[5]&r_0_addr[11],
r_2_addr[13]&r_1_addr[5]&r_0_addr[10],
r_2_addr[13]&r_1_addr[5]&r_0_addr[9],
r_2_addr[13]&r_1_addr[5]&r_0_addr[8],
r_2_addr[13]&r_1_addr[5]&r_0_addr[7],
r_2_addr[13]&r_1_addr[5]&r_0_addr[6],
r_2_addr[13]&r_1_addr[5]&r_0_addr[5],
r_2_addr[13]&r_1_addr[5]&r_0_addr[4],
r_2_addr[13]&r_1_addr[5]&r_0_addr[3],
r_2_addr[13]&r_1_addr[5]&r_0_addr[2],
r_2_addr[13]&r_1_addr[5]&r_0_addr[1],
r_2_addr[13]&r_1_addr[5]&r_0_addr[0],
r_2_addr[13]&r_1_addr[4]&r_0_addr[15],
r_2_addr[13]&r_1_addr[4]&r_0_addr[14],
r_2_addr[13]&r_1_addr[4]&r_0_addr[13],
r_2_addr[13]&r_1_addr[4]&r_0_addr[12],
r_2_addr[13]&r_1_addr[4]&r_0_addr[11],
r_2_addr[13]&r_1_addr[4]&r_0_addr[10],
r_2_addr[13]&r_1_addr[4]&r_0_addr[9],
r_2_addr[13]&r_1_addr[4]&r_0_addr[8],
r_2_addr[13]&r_1_addr[4]&r_0_addr[7],
r_2_addr[13]&r_1_addr[4]&r_0_addr[6],
r_2_addr[13]&r_1_addr[4]&r_0_addr[5],
r_2_addr[13]&r_1_addr[4]&r_0_addr[4],
r_2_addr[13]&r_1_addr[4]&r_0_addr[3],
r_2_addr[13]&r_1_addr[4]&r_0_addr[2],
r_2_addr[13]&r_1_addr[4]&r_0_addr[1],
r_2_addr[13]&r_1_addr[4]&r_0_addr[0],
r_2_addr[13]&r_1_addr[3]&r_0_addr[15],
r_2_addr[13]&r_1_addr[3]&r_0_addr[14],
r_2_addr[13]&r_1_addr[3]&r_0_addr[13],
r_2_addr[13]&r_1_addr[3]&r_0_addr[12],
r_2_addr[13]&r_1_addr[3]&r_0_addr[11],
r_2_addr[13]&r_1_addr[3]&r_0_addr[10],
r_2_addr[13]&r_1_addr[3]&r_0_addr[9],
r_2_addr[13]&r_1_addr[3]&r_0_addr[8],
r_2_addr[13]&r_1_addr[3]&r_0_addr[7],
r_2_addr[13]&r_1_addr[3]&r_0_addr[6],
r_2_addr[13]&r_1_addr[3]&r_0_addr[5],
r_2_addr[13]&r_1_addr[3]&r_0_addr[4],
r_2_addr[13]&r_1_addr[3]&r_0_addr[3],
r_2_addr[13]&r_1_addr[3]&r_0_addr[2],
r_2_addr[13]&r_1_addr[3]&r_0_addr[1],
r_2_addr[13]&r_1_addr[3]&r_0_addr[0],
r_2_addr[13]&r_1_addr[2]&r_0_addr[15],
r_2_addr[13]&r_1_addr[2]&r_0_addr[14],
r_2_addr[13]&r_1_addr[2]&r_0_addr[13],
r_2_addr[13]&r_1_addr[2]&r_0_addr[12],
r_2_addr[13]&r_1_addr[2]&r_0_addr[11],
r_2_addr[13]&r_1_addr[2]&r_0_addr[10],
r_2_addr[13]&r_1_addr[2]&r_0_addr[9],
r_2_addr[13]&r_1_addr[2]&r_0_addr[8],
r_2_addr[13]&r_1_addr[2]&r_0_addr[7],
r_2_addr[13]&r_1_addr[2]&r_0_addr[6],
r_2_addr[13]&r_1_addr[2]&r_0_addr[5],
r_2_addr[13]&r_1_addr[2]&r_0_addr[4],
r_2_addr[13]&r_1_addr[2]&r_0_addr[3],
r_2_addr[13]&r_1_addr[2]&r_0_addr[2],
r_2_addr[13]&r_1_addr[2]&r_0_addr[1],
r_2_addr[13]&r_1_addr[2]&r_0_addr[0],
r_2_addr[13]&r_1_addr[1]&r_0_addr[15],
r_2_addr[13]&r_1_addr[1]&r_0_addr[14],
r_2_addr[13]&r_1_addr[1]&r_0_addr[13],
r_2_addr[13]&r_1_addr[1]&r_0_addr[12],
r_2_addr[13]&r_1_addr[1]&r_0_addr[11],
r_2_addr[13]&r_1_addr[1]&r_0_addr[10],
r_2_addr[13]&r_1_addr[1]&r_0_addr[9],
r_2_addr[13]&r_1_addr[1]&r_0_addr[8],
r_2_addr[13]&r_1_addr[1]&r_0_addr[7],
r_2_addr[13]&r_1_addr[1]&r_0_addr[6],
r_2_addr[13]&r_1_addr[1]&r_0_addr[5],
r_2_addr[13]&r_1_addr[1]&r_0_addr[4],
r_2_addr[13]&r_1_addr[1]&r_0_addr[3],
r_2_addr[13]&r_1_addr[1]&r_0_addr[2],
r_2_addr[13]&r_1_addr[1]&r_0_addr[1],
r_2_addr[13]&r_1_addr[1]&r_0_addr[0],
r_2_addr[13]&r_1_addr[0]&r_0_addr[15],
r_2_addr[13]&r_1_addr[0]&r_0_addr[14],
r_2_addr[13]&r_1_addr[0]&r_0_addr[13],
r_2_addr[13]&r_1_addr[0]&r_0_addr[12],
r_2_addr[13]&r_1_addr[0]&r_0_addr[11],
r_2_addr[13]&r_1_addr[0]&r_0_addr[10],
r_2_addr[13]&r_1_addr[0]&r_0_addr[9],
r_2_addr[13]&r_1_addr[0]&r_0_addr[8],
r_2_addr[13]&r_1_addr[0]&r_0_addr[7],
r_2_addr[13]&r_1_addr[0]&r_0_addr[6],
r_2_addr[13]&r_1_addr[0]&r_0_addr[5],
r_2_addr[13]&r_1_addr[0]&r_0_addr[4],
r_2_addr[13]&r_1_addr[0]&r_0_addr[3],
r_2_addr[13]&r_1_addr[0]&r_0_addr[2],
r_2_addr[13]&r_1_addr[0]&r_0_addr[1],
r_2_addr[13]&r_1_addr[0]&r_0_addr[0],
r_2_addr[12]&r_1_addr[15]&r_0_addr[15],
r_2_addr[12]&r_1_addr[15]&r_0_addr[14],
r_2_addr[12]&r_1_addr[15]&r_0_addr[13],
r_2_addr[12]&r_1_addr[15]&r_0_addr[12],
r_2_addr[12]&r_1_addr[15]&r_0_addr[11],
r_2_addr[12]&r_1_addr[15]&r_0_addr[10],
r_2_addr[12]&r_1_addr[15]&r_0_addr[9],
r_2_addr[12]&r_1_addr[15]&r_0_addr[8],
r_2_addr[12]&r_1_addr[15]&r_0_addr[7],
r_2_addr[12]&r_1_addr[15]&r_0_addr[6],
r_2_addr[12]&r_1_addr[15]&r_0_addr[5],
r_2_addr[12]&r_1_addr[15]&r_0_addr[4],
r_2_addr[12]&r_1_addr[15]&r_0_addr[3],
r_2_addr[12]&r_1_addr[15]&r_0_addr[2],
r_2_addr[12]&r_1_addr[15]&r_0_addr[1],
r_2_addr[12]&r_1_addr[15]&r_0_addr[0],
r_2_addr[12]&r_1_addr[14]&r_0_addr[15],
r_2_addr[12]&r_1_addr[14]&r_0_addr[14],
r_2_addr[12]&r_1_addr[14]&r_0_addr[13],
r_2_addr[12]&r_1_addr[14]&r_0_addr[12],
r_2_addr[12]&r_1_addr[14]&r_0_addr[11],
r_2_addr[12]&r_1_addr[14]&r_0_addr[10],
r_2_addr[12]&r_1_addr[14]&r_0_addr[9],
r_2_addr[12]&r_1_addr[14]&r_0_addr[8],
r_2_addr[12]&r_1_addr[14]&r_0_addr[7],
r_2_addr[12]&r_1_addr[14]&r_0_addr[6],
r_2_addr[12]&r_1_addr[14]&r_0_addr[5],
r_2_addr[12]&r_1_addr[14]&r_0_addr[4],
r_2_addr[12]&r_1_addr[14]&r_0_addr[3],
r_2_addr[12]&r_1_addr[14]&r_0_addr[2],
r_2_addr[12]&r_1_addr[14]&r_0_addr[1],
r_2_addr[12]&r_1_addr[14]&r_0_addr[0],
r_2_addr[12]&r_1_addr[13]&r_0_addr[15],
r_2_addr[12]&r_1_addr[13]&r_0_addr[14],
r_2_addr[12]&r_1_addr[13]&r_0_addr[13],
r_2_addr[12]&r_1_addr[13]&r_0_addr[12],
r_2_addr[12]&r_1_addr[13]&r_0_addr[11],
r_2_addr[12]&r_1_addr[13]&r_0_addr[10],
r_2_addr[12]&r_1_addr[13]&r_0_addr[9],
r_2_addr[12]&r_1_addr[13]&r_0_addr[8],
r_2_addr[12]&r_1_addr[13]&r_0_addr[7],
r_2_addr[12]&r_1_addr[13]&r_0_addr[6],
r_2_addr[12]&r_1_addr[13]&r_0_addr[5],
r_2_addr[12]&r_1_addr[13]&r_0_addr[4],
r_2_addr[12]&r_1_addr[13]&r_0_addr[3],
r_2_addr[12]&r_1_addr[13]&r_0_addr[2],
r_2_addr[12]&r_1_addr[13]&r_0_addr[1],
r_2_addr[12]&r_1_addr[13]&r_0_addr[0],
r_2_addr[12]&r_1_addr[12]&r_0_addr[15],
r_2_addr[12]&r_1_addr[12]&r_0_addr[14],
r_2_addr[12]&r_1_addr[12]&r_0_addr[13],
r_2_addr[12]&r_1_addr[12]&r_0_addr[12],
r_2_addr[12]&r_1_addr[12]&r_0_addr[11],
r_2_addr[12]&r_1_addr[12]&r_0_addr[10],
r_2_addr[12]&r_1_addr[12]&r_0_addr[9],
r_2_addr[12]&r_1_addr[12]&r_0_addr[8],
r_2_addr[12]&r_1_addr[12]&r_0_addr[7],
r_2_addr[12]&r_1_addr[12]&r_0_addr[6],
r_2_addr[12]&r_1_addr[12]&r_0_addr[5],
r_2_addr[12]&r_1_addr[12]&r_0_addr[4],
r_2_addr[12]&r_1_addr[12]&r_0_addr[3],
r_2_addr[12]&r_1_addr[12]&r_0_addr[2],
r_2_addr[12]&r_1_addr[12]&r_0_addr[1],
r_2_addr[12]&r_1_addr[12]&r_0_addr[0],
r_2_addr[12]&r_1_addr[11]&r_0_addr[15],
r_2_addr[12]&r_1_addr[11]&r_0_addr[14],
r_2_addr[12]&r_1_addr[11]&r_0_addr[13],
r_2_addr[12]&r_1_addr[11]&r_0_addr[12],
r_2_addr[12]&r_1_addr[11]&r_0_addr[11],
r_2_addr[12]&r_1_addr[11]&r_0_addr[10],
r_2_addr[12]&r_1_addr[11]&r_0_addr[9],
r_2_addr[12]&r_1_addr[11]&r_0_addr[8],
r_2_addr[12]&r_1_addr[11]&r_0_addr[7],
r_2_addr[12]&r_1_addr[11]&r_0_addr[6],
r_2_addr[12]&r_1_addr[11]&r_0_addr[5],
r_2_addr[12]&r_1_addr[11]&r_0_addr[4],
r_2_addr[12]&r_1_addr[11]&r_0_addr[3],
r_2_addr[12]&r_1_addr[11]&r_0_addr[2],
r_2_addr[12]&r_1_addr[11]&r_0_addr[1],
r_2_addr[12]&r_1_addr[11]&r_0_addr[0],
r_2_addr[12]&r_1_addr[10]&r_0_addr[15],
r_2_addr[12]&r_1_addr[10]&r_0_addr[14],
r_2_addr[12]&r_1_addr[10]&r_0_addr[13],
r_2_addr[12]&r_1_addr[10]&r_0_addr[12],
r_2_addr[12]&r_1_addr[10]&r_0_addr[11],
r_2_addr[12]&r_1_addr[10]&r_0_addr[10],
r_2_addr[12]&r_1_addr[10]&r_0_addr[9],
r_2_addr[12]&r_1_addr[10]&r_0_addr[8],
r_2_addr[12]&r_1_addr[10]&r_0_addr[7],
r_2_addr[12]&r_1_addr[10]&r_0_addr[6],
r_2_addr[12]&r_1_addr[10]&r_0_addr[5],
r_2_addr[12]&r_1_addr[10]&r_0_addr[4],
r_2_addr[12]&r_1_addr[10]&r_0_addr[3],
r_2_addr[12]&r_1_addr[10]&r_0_addr[2],
r_2_addr[12]&r_1_addr[10]&r_0_addr[1],
r_2_addr[12]&r_1_addr[10]&r_0_addr[0],
r_2_addr[12]&r_1_addr[9]&r_0_addr[15],
r_2_addr[12]&r_1_addr[9]&r_0_addr[14],
r_2_addr[12]&r_1_addr[9]&r_0_addr[13],
r_2_addr[12]&r_1_addr[9]&r_0_addr[12],
r_2_addr[12]&r_1_addr[9]&r_0_addr[11],
r_2_addr[12]&r_1_addr[9]&r_0_addr[10],
r_2_addr[12]&r_1_addr[9]&r_0_addr[9],
r_2_addr[12]&r_1_addr[9]&r_0_addr[8],
r_2_addr[12]&r_1_addr[9]&r_0_addr[7],
r_2_addr[12]&r_1_addr[9]&r_0_addr[6],
r_2_addr[12]&r_1_addr[9]&r_0_addr[5],
r_2_addr[12]&r_1_addr[9]&r_0_addr[4],
r_2_addr[12]&r_1_addr[9]&r_0_addr[3],
r_2_addr[12]&r_1_addr[9]&r_0_addr[2],
r_2_addr[12]&r_1_addr[9]&r_0_addr[1],
r_2_addr[12]&r_1_addr[9]&r_0_addr[0],
r_2_addr[12]&r_1_addr[8]&r_0_addr[15],
r_2_addr[12]&r_1_addr[8]&r_0_addr[14],
r_2_addr[12]&r_1_addr[8]&r_0_addr[13],
r_2_addr[12]&r_1_addr[8]&r_0_addr[12],
r_2_addr[12]&r_1_addr[8]&r_0_addr[11],
r_2_addr[12]&r_1_addr[8]&r_0_addr[10],
r_2_addr[12]&r_1_addr[8]&r_0_addr[9],
r_2_addr[12]&r_1_addr[8]&r_0_addr[8],
r_2_addr[12]&r_1_addr[8]&r_0_addr[7],
r_2_addr[12]&r_1_addr[8]&r_0_addr[6],
r_2_addr[12]&r_1_addr[8]&r_0_addr[5],
r_2_addr[12]&r_1_addr[8]&r_0_addr[4],
r_2_addr[12]&r_1_addr[8]&r_0_addr[3],
r_2_addr[12]&r_1_addr[8]&r_0_addr[2],
r_2_addr[12]&r_1_addr[8]&r_0_addr[1],
r_2_addr[12]&r_1_addr[8]&r_0_addr[0],
r_2_addr[12]&r_1_addr[7]&r_0_addr[15],
r_2_addr[12]&r_1_addr[7]&r_0_addr[14],
r_2_addr[12]&r_1_addr[7]&r_0_addr[13],
r_2_addr[12]&r_1_addr[7]&r_0_addr[12],
r_2_addr[12]&r_1_addr[7]&r_0_addr[11],
r_2_addr[12]&r_1_addr[7]&r_0_addr[10],
r_2_addr[12]&r_1_addr[7]&r_0_addr[9],
r_2_addr[12]&r_1_addr[7]&r_0_addr[8],
r_2_addr[12]&r_1_addr[7]&r_0_addr[7],
r_2_addr[12]&r_1_addr[7]&r_0_addr[6],
r_2_addr[12]&r_1_addr[7]&r_0_addr[5],
r_2_addr[12]&r_1_addr[7]&r_0_addr[4],
r_2_addr[12]&r_1_addr[7]&r_0_addr[3],
r_2_addr[12]&r_1_addr[7]&r_0_addr[2],
r_2_addr[12]&r_1_addr[7]&r_0_addr[1],
r_2_addr[12]&r_1_addr[7]&r_0_addr[0],
r_2_addr[12]&r_1_addr[6]&r_0_addr[15],
r_2_addr[12]&r_1_addr[6]&r_0_addr[14],
r_2_addr[12]&r_1_addr[6]&r_0_addr[13],
r_2_addr[12]&r_1_addr[6]&r_0_addr[12],
r_2_addr[12]&r_1_addr[6]&r_0_addr[11],
r_2_addr[12]&r_1_addr[6]&r_0_addr[10],
r_2_addr[12]&r_1_addr[6]&r_0_addr[9],
r_2_addr[12]&r_1_addr[6]&r_0_addr[8],
r_2_addr[12]&r_1_addr[6]&r_0_addr[7],
r_2_addr[12]&r_1_addr[6]&r_0_addr[6],
r_2_addr[12]&r_1_addr[6]&r_0_addr[5],
r_2_addr[12]&r_1_addr[6]&r_0_addr[4],
r_2_addr[12]&r_1_addr[6]&r_0_addr[3],
r_2_addr[12]&r_1_addr[6]&r_0_addr[2],
r_2_addr[12]&r_1_addr[6]&r_0_addr[1],
r_2_addr[12]&r_1_addr[6]&r_0_addr[0],
r_2_addr[12]&r_1_addr[5]&r_0_addr[15],
r_2_addr[12]&r_1_addr[5]&r_0_addr[14],
r_2_addr[12]&r_1_addr[5]&r_0_addr[13],
r_2_addr[12]&r_1_addr[5]&r_0_addr[12],
r_2_addr[12]&r_1_addr[5]&r_0_addr[11],
r_2_addr[12]&r_1_addr[5]&r_0_addr[10],
r_2_addr[12]&r_1_addr[5]&r_0_addr[9],
r_2_addr[12]&r_1_addr[5]&r_0_addr[8],
r_2_addr[12]&r_1_addr[5]&r_0_addr[7],
r_2_addr[12]&r_1_addr[5]&r_0_addr[6],
r_2_addr[12]&r_1_addr[5]&r_0_addr[5],
r_2_addr[12]&r_1_addr[5]&r_0_addr[4],
r_2_addr[12]&r_1_addr[5]&r_0_addr[3],
r_2_addr[12]&r_1_addr[5]&r_0_addr[2],
r_2_addr[12]&r_1_addr[5]&r_0_addr[1],
r_2_addr[12]&r_1_addr[5]&r_0_addr[0],
r_2_addr[12]&r_1_addr[4]&r_0_addr[15],
r_2_addr[12]&r_1_addr[4]&r_0_addr[14],
r_2_addr[12]&r_1_addr[4]&r_0_addr[13],
r_2_addr[12]&r_1_addr[4]&r_0_addr[12],
r_2_addr[12]&r_1_addr[4]&r_0_addr[11],
r_2_addr[12]&r_1_addr[4]&r_0_addr[10],
r_2_addr[12]&r_1_addr[4]&r_0_addr[9],
r_2_addr[12]&r_1_addr[4]&r_0_addr[8],
r_2_addr[12]&r_1_addr[4]&r_0_addr[7],
r_2_addr[12]&r_1_addr[4]&r_0_addr[6],
r_2_addr[12]&r_1_addr[4]&r_0_addr[5],
r_2_addr[12]&r_1_addr[4]&r_0_addr[4],
r_2_addr[12]&r_1_addr[4]&r_0_addr[3],
r_2_addr[12]&r_1_addr[4]&r_0_addr[2],
r_2_addr[12]&r_1_addr[4]&r_0_addr[1],
r_2_addr[12]&r_1_addr[4]&r_0_addr[0],
r_2_addr[12]&r_1_addr[3]&r_0_addr[15],
r_2_addr[12]&r_1_addr[3]&r_0_addr[14],
r_2_addr[12]&r_1_addr[3]&r_0_addr[13],
r_2_addr[12]&r_1_addr[3]&r_0_addr[12],
r_2_addr[12]&r_1_addr[3]&r_0_addr[11],
r_2_addr[12]&r_1_addr[3]&r_0_addr[10],
r_2_addr[12]&r_1_addr[3]&r_0_addr[9],
r_2_addr[12]&r_1_addr[3]&r_0_addr[8],
r_2_addr[12]&r_1_addr[3]&r_0_addr[7],
r_2_addr[12]&r_1_addr[3]&r_0_addr[6],
r_2_addr[12]&r_1_addr[3]&r_0_addr[5],
r_2_addr[12]&r_1_addr[3]&r_0_addr[4],
r_2_addr[12]&r_1_addr[3]&r_0_addr[3],
r_2_addr[12]&r_1_addr[3]&r_0_addr[2],
r_2_addr[12]&r_1_addr[3]&r_0_addr[1],
r_2_addr[12]&r_1_addr[3]&r_0_addr[0],
r_2_addr[12]&r_1_addr[2]&r_0_addr[15],
r_2_addr[12]&r_1_addr[2]&r_0_addr[14],
r_2_addr[12]&r_1_addr[2]&r_0_addr[13],
r_2_addr[12]&r_1_addr[2]&r_0_addr[12],
r_2_addr[12]&r_1_addr[2]&r_0_addr[11],
r_2_addr[12]&r_1_addr[2]&r_0_addr[10],
r_2_addr[12]&r_1_addr[2]&r_0_addr[9],
r_2_addr[12]&r_1_addr[2]&r_0_addr[8],
r_2_addr[12]&r_1_addr[2]&r_0_addr[7],
r_2_addr[12]&r_1_addr[2]&r_0_addr[6],
r_2_addr[12]&r_1_addr[2]&r_0_addr[5],
r_2_addr[12]&r_1_addr[2]&r_0_addr[4],
r_2_addr[12]&r_1_addr[2]&r_0_addr[3],
r_2_addr[12]&r_1_addr[2]&r_0_addr[2],
r_2_addr[12]&r_1_addr[2]&r_0_addr[1],
r_2_addr[12]&r_1_addr[2]&r_0_addr[0],
r_2_addr[12]&r_1_addr[1]&r_0_addr[15],
r_2_addr[12]&r_1_addr[1]&r_0_addr[14],
r_2_addr[12]&r_1_addr[1]&r_0_addr[13],
r_2_addr[12]&r_1_addr[1]&r_0_addr[12],
r_2_addr[12]&r_1_addr[1]&r_0_addr[11],
r_2_addr[12]&r_1_addr[1]&r_0_addr[10],
r_2_addr[12]&r_1_addr[1]&r_0_addr[9],
r_2_addr[12]&r_1_addr[1]&r_0_addr[8],
r_2_addr[12]&r_1_addr[1]&r_0_addr[7],
r_2_addr[12]&r_1_addr[1]&r_0_addr[6],
r_2_addr[12]&r_1_addr[1]&r_0_addr[5],
r_2_addr[12]&r_1_addr[1]&r_0_addr[4],
r_2_addr[12]&r_1_addr[1]&r_0_addr[3],
r_2_addr[12]&r_1_addr[1]&r_0_addr[2],
r_2_addr[12]&r_1_addr[1]&r_0_addr[1],
r_2_addr[12]&r_1_addr[1]&r_0_addr[0],
r_2_addr[12]&r_1_addr[0]&r_0_addr[15],
r_2_addr[12]&r_1_addr[0]&r_0_addr[14],
r_2_addr[12]&r_1_addr[0]&r_0_addr[13],
r_2_addr[12]&r_1_addr[0]&r_0_addr[12],
r_2_addr[12]&r_1_addr[0]&r_0_addr[11],
r_2_addr[12]&r_1_addr[0]&r_0_addr[10],
r_2_addr[12]&r_1_addr[0]&r_0_addr[9],
r_2_addr[12]&r_1_addr[0]&r_0_addr[8],
r_2_addr[12]&r_1_addr[0]&r_0_addr[7],
r_2_addr[12]&r_1_addr[0]&r_0_addr[6],
r_2_addr[12]&r_1_addr[0]&r_0_addr[5],
r_2_addr[12]&r_1_addr[0]&r_0_addr[4],
r_2_addr[12]&r_1_addr[0]&r_0_addr[3],
r_2_addr[12]&r_1_addr[0]&r_0_addr[2],
r_2_addr[12]&r_1_addr[0]&r_0_addr[1],
r_2_addr[12]&r_1_addr[0]&r_0_addr[0],
r_2_addr[11]&r_1_addr[15]&r_0_addr[15],
r_2_addr[11]&r_1_addr[15]&r_0_addr[14],
r_2_addr[11]&r_1_addr[15]&r_0_addr[13],
r_2_addr[11]&r_1_addr[15]&r_0_addr[12],
r_2_addr[11]&r_1_addr[15]&r_0_addr[11],
r_2_addr[11]&r_1_addr[15]&r_0_addr[10],
r_2_addr[11]&r_1_addr[15]&r_0_addr[9],
r_2_addr[11]&r_1_addr[15]&r_0_addr[8],
r_2_addr[11]&r_1_addr[15]&r_0_addr[7],
r_2_addr[11]&r_1_addr[15]&r_0_addr[6],
r_2_addr[11]&r_1_addr[15]&r_0_addr[5],
r_2_addr[11]&r_1_addr[15]&r_0_addr[4],
r_2_addr[11]&r_1_addr[15]&r_0_addr[3],
r_2_addr[11]&r_1_addr[15]&r_0_addr[2],
r_2_addr[11]&r_1_addr[15]&r_0_addr[1],
r_2_addr[11]&r_1_addr[15]&r_0_addr[0],
r_2_addr[11]&r_1_addr[14]&r_0_addr[15],
r_2_addr[11]&r_1_addr[14]&r_0_addr[14],
r_2_addr[11]&r_1_addr[14]&r_0_addr[13],
r_2_addr[11]&r_1_addr[14]&r_0_addr[12],
r_2_addr[11]&r_1_addr[14]&r_0_addr[11],
r_2_addr[11]&r_1_addr[14]&r_0_addr[10],
r_2_addr[11]&r_1_addr[14]&r_0_addr[9],
r_2_addr[11]&r_1_addr[14]&r_0_addr[8],
r_2_addr[11]&r_1_addr[14]&r_0_addr[7],
r_2_addr[11]&r_1_addr[14]&r_0_addr[6],
r_2_addr[11]&r_1_addr[14]&r_0_addr[5],
r_2_addr[11]&r_1_addr[14]&r_0_addr[4],
r_2_addr[11]&r_1_addr[14]&r_0_addr[3],
r_2_addr[11]&r_1_addr[14]&r_0_addr[2],
r_2_addr[11]&r_1_addr[14]&r_0_addr[1],
r_2_addr[11]&r_1_addr[14]&r_0_addr[0],
r_2_addr[11]&r_1_addr[13]&r_0_addr[15],
r_2_addr[11]&r_1_addr[13]&r_0_addr[14],
r_2_addr[11]&r_1_addr[13]&r_0_addr[13],
r_2_addr[11]&r_1_addr[13]&r_0_addr[12],
r_2_addr[11]&r_1_addr[13]&r_0_addr[11],
r_2_addr[11]&r_1_addr[13]&r_0_addr[10],
r_2_addr[11]&r_1_addr[13]&r_0_addr[9],
r_2_addr[11]&r_1_addr[13]&r_0_addr[8],
r_2_addr[11]&r_1_addr[13]&r_0_addr[7],
r_2_addr[11]&r_1_addr[13]&r_0_addr[6],
r_2_addr[11]&r_1_addr[13]&r_0_addr[5],
r_2_addr[11]&r_1_addr[13]&r_0_addr[4],
r_2_addr[11]&r_1_addr[13]&r_0_addr[3],
r_2_addr[11]&r_1_addr[13]&r_0_addr[2],
r_2_addr[11]&r_1_addr[13]&r_0_addr[1],
r_2_addr[11]&r_1_addr[13]&r_0_addr[0],
r_2_addr[11]&r_1_addr[12]&r_0_addr[15],
r_2_addr[11]&r_1_addr[12]&r_0_addr[14],
r_2_addr[11]&r_1_addr[12]&r_0_addr[13],
r_2_addr[11]&r_1_addr[12]&r_0_addr[12],
r_2_addr[11]&r_1_addr[12]&r_0_addr[11],
r_2_addr[11]&r_1_addr[12]&r_0_addr[10],
r_2_addr[11]&r_1_addr[12]&r_0_addr[9],
r_2_addr[11]&r_1_addr[12]&r_0_addr[8],
r_2_addr[11]&r_1_addr[12]&r_0_addr[7],
r_2_addr[11]&r_1_addr[12]&r_0_addr[6],
r_2_addr[11]&r_1_addr[12]&r_0_addr[5],
r_2_addr[11]&r_1_addr[12]&r_0_addr[4],
r_2_addr[11]&r_1_addr[12]&r_0_addr[3],
r_2_addr[11]&r_1_addr[12]&r_0_addr[2],
r_2_addr[11]&r_1_addr[12]&r_0_addr[1],
r_2_addr[11]&r_1_addr[12]&r_0_addr[0],
r_2_addr[11]&r_1_addr[11]&r_0_addr[15],
r_2_addr[11]&r_1_addr[11]&r_0_addr[14],
r_2_addr[11]&r_1_addr[11]&r_0_addr[13],
r_2_addr[11]&r_1_addr[11]&r_0_addr[12],
r_2_addr[11]&r_1_addr[11]&r_0_addr[11],
r_2_addr[11]&r_1_addr[11]&r_0_addr[10],
r_2_addr[11]&r_1_addr[11]&r_0_addr[9],
r_2_addr[11]&r_1_addr[11]&r_0_addr[8],
r_2_addr[11]&r_1_addr[11]&r_0_addr[7],
r_2_addr[11]&r_1_addr[11]&r_0_addr[6],
r_2_addr[11]&r_1_addr[11]&r_0_addr[5],
r_2_addr[11]&r_1_addr[11]&r_0_addr[4],
r_2_addr[11]&r_1_addr[11]&r_0_addr[3],
r_2_addr[11]&r_1_addr[11]&r_0_addr[2],
r_2_addr[11]&r_1_addr[11]&r_0_addr[1],
r_2_addr[11]&r_1_addr[11]&r_0_addr[0],
r_2_addr[11]&r_1_addr[10]&r_0_addr[15],
r_2_addr[11]&r_1_addr[10]&r_0_addr[14],
r_2_addr[11]&r_1_addr[10]&r_0_addr[13],
r_2_addr[11]&r_1_addr[10]&r_0_addr[12],
r_2_addr[11]&r_1_addr[10]&r_0_addr[11],
r_2_addr[11]&r_1_addr[10]&r_0_addr[10],
r_2_addr[11]&r_1_addr[10]&r_0_addr[9],
r_2_addr[11]&r_1_addr[10]&r_0_addr[8],
r_2_addr[11]&r_1_addr[10]&r_0_addr[7],
r_2_addr[11]&r_1_addr[10]&r_0_addr[6],
r_2_addr[11]&r_1_addr[10]&r_0_addr[5],
r_2_addr[11]&r_1_addr[10]&r_0_addr[4],
r_2_addr[11]&r_1_addr[10]&r_0_addr[3],
r_2_addr[11]&r_1_addr[10]&r_0_addr[2],
r_2_addr[11]&r_1_addr[10]&r_0_addr[1],
r_2_addr[11]&r_1_addr[10]&r_0_addr[0],
r_2_addr[11]&r_1_addr[9]&r_0_addr[15],
r_2_addr[11]&r_1_addr[9]&r_0_addr[14],
r_2_addr[11]&r_1_addr[9]&r_0_addr[13],
r_2_addr[11]&r_1_addr[9]&r_0_addr[12],
r_2_addr[11]&r_1_addr[9]&r_0_addr[11],
r_2_addr[11]&r_1_addr[9]&r_0_addr[10],
r_2_addr[11]&r_1_addr[9]&r_0_addr[9],
r_2_addr[11]&r_1_addr[9]&r_0_addr[8],
r_2_addr[11]&r_1_addr[9]&r_0_addr[7],
r_2_addr[11]&r_1_addr[9]&r_0_addr[6],
r_2_addr[11]&r_1_addr[9]&r_0_addr[5],
r_2_addr[11]&r_1_addr[9]&r_0_addr[4],
r_2_addr[11]&r_1_addr[9]&r_0_addr[3],
r_2_addr[11]&r_1_addr[9]&r_0_addr[2],
r_2_addr[11]&r_1_addr[9]&r_0_addr[1],
r_2_addr[11]&r_1_addr[9]&r_0_addr[0],
r_2_addr[11]&r_1_addr[8]&r_0_addr[15],
r_2_addr[11]&r_1_addr[8]&r_0_addr[14],
r_2_addr[11]&r_1_addr[8]&r_0_addr[13],
r_2_addr[11]&r_1_addr[8]&r_0_addr[12],
r_2_addr[11]&r_1_addr[8]&r_0_addr[11],
r_2_addr[11]&r_1_addr[8]&r_0_addr[10],
r_2_addr[11]&r_1_addr[8]&r_0_addr[9],
r_2_addr[11]&r_1_addr[8]&r_0_addr[8],
r_2_addr[11]&r_1_addr[8]&r_0_addr[7],
r_2_addr[11]&r_1_addr[8]&r_0_addr[6],
r_2_addr[11]&r_1_addr[8]&r_0_addr[5],
r_2_addr[11]&r_1_addr[8]&r_0_addr[4],
r_2_addr[11]&r_1_addr[8]&r_0_addr[3],
r_2_addr[11]&r_1_addr[8]&r_0_addr[2],
r_2_addr[11]&r_1_addr[8]&r_0_addr[1],
r_2_addr[11]&r_1_addr[8]&r_0_addr[0],
r_2_addr[11]&r_1_addr[7]&r_0_addr[15],
r_2_addr[11]&r_1_addr[7]&r_0_addr[14],
r_2_addr[11]&r_1_addr[7]&r_0_addr[13],
r_2_addr[11]&r_1_addr[7]&r_0_addr[12],
r_2_addr[11]&r_1_addr[7]&r_0_addr[11],
r_2_addr[11]&r_1_addr[7]&r_0_addr[10],
r_2_addr[11]&r_1_addr[7]&r_0_addr[9],
r_2_addr[11]&r_1_addr[7]&r_0_addr[8],
r_2_addr[11]&r_1_addr[7]&r_0_addr[7],
r_2_addr[11]&r_1_addr[7]&r_0_addr[6],
r_2_addr[11]&r_1_addr[7]&r_0_addr[5],
r_2_addr[11]&r_1_addr[7]&r_0_addr[4],
r_2_addr[11]&r_1_addr[7]&r_0_addr[3],
r_2_addr[11]&r_1_addr[7]&r_0_addr[2],
r_2_addr[11]&r_1_addr[7]&r_0_addr[1],
r_2_addr[11]&r_1_addr[7]&r_0_addr[0],
r_2_addr[11]&r_1_addr[6]&r_0_addr[15],
r_2_addr[11]&r_1_addr[6]&r_0_addr[14],
r_2_addr[11]&r_1_addr[6]&r_0_addr[13],
r_2_addr[11]&r_1_addr[6]&r_0_addr[12],
r_2_addr[11]&r_1_addr[6]&r_0_addr[11],
r_2_addr[11]&r_1_addr[6]&r_0_addr[10],
r_2_addr[11]&r_1_addr[6]&r_0_addr[9],
r_2_addr[11]&r_1_addr[6]&r_0_addr[8],
r_2_addr[11]&r_1_addr[6]&r_0_addr[7],
r_2_addr[11]&r_1_addr[6]&r_0_addr[6],
r_2_addr[11]&r_1_addr[6]&r_0_addr[5],
r_2_addr[11]&r_1_addr[6]&r_0_addr[4],
r_2_addr[11]&r_1_addr[6]&r_0_addr[3],
r_2_addr[11]&r_1_addr[6]&r_0_addr[2],
r_2_addr[11]&r_1_addr[6]&r_0_addr[1],
r_2_addr[11]&r_1_addr[6]&r_0_addr[0],
r_2_addr[11]&r_1_addr[5]&r_0_addr[15],
r_2_addr[11]&r_1_addr[5]&r_0_addr[14],
r_2_addr[11]&r_1_addr[5]&r_0_addr[13],
r_2_addr[11]&r_1_addr[5]&r_0_addr[12],
r_2_addr[11]&r_1_addr[5]&r_0_addr[11],
r_2_addr[11]&r_1_addr[5]&r_0_addr[10],
r_2_addr[11]&r_1_addr[5]&r_0_addr[9],
r_2_addr[11]&r_1_addr[5]&r_0_addr[8],
r_2_addr[11]&r_1_addr[5]&r_0_addr[7],
r_2_addr[11]&r_1_addr[5]&r_0_addr[6],
r_2_addr[11]&r_1_addr[5]&r_0_addr[5],
r_2_addr[11]&r_1_addr[5]&r_0_addr[4],
r_2_addr[11]&r_1_addr[5]&r_0_addr[3],
r_2_addr[11]&r_1_addr[5]&r_0_addr[2],
r_2_addr[11]&r_1_addr[5]&r_0_addr[1],
r_2_addr[11]&r_1_addr[5]&r_0_addr[0],
r_2_addr[11]&r_1_addr[4]&r_0_addr[15],
r_2_addr[11]&r_1_addr[4]&r_0_addr[14],
r_2_addr[11]&r_1_addr[4]&r_0_addr[13],
r_2_addr[11]&r_1_addr[4]&r_0_addr[12],
r_2_addr[11]&r_1_addr[4]&r_0_addr[11],
r_2_addr[11]&r_1_addr[4]&r_0_addr[10],
r_2_addr[11]&r_1_addr[4]&r_0_addr[9],
r_2_addr[11]&r_1_addr[4]&r_0_addr[8],
r_2_addr[11]&r_1_addr[4]&r_0_addr[7],
r_2_addr[11]&r_1_addr[4]&r_0_addr[6],
r_2_addr[11]&r_1_addr[4]&r_0_addr[5],
r_2_addr[11]&r_1_addr[4]&r_0_addr[4],
r_2_addr[11]&r_1_addr[4]&r_0_addr[3],
r_2_addr[11]&r_1_addr[4]&r_0_addr[2],
r_2_addr[11]&r_1_addr[4]&r_0_addr[1],
r_2_addr[11]&r_1_addr[4]&r_0_addr[0],
r_2_addr[11]&r_1_addr[3]&r_0_addr[15],
r_2_addr[11]&r_1_addr[3]&r_0_addr[14],
r_2_addr[11]&r_1_addr[3]&r_0_addr[13],
r_2_addr[11]&r_1_addr[3]&r_0_addr[12],
r_2_addr[11]&r_1_addr[3]&r_0_addr[11],
r_2_addr[11]&r_1_addr[3]&r_0_addr[10],
r_2_addr[11]&r_1_addr[3]&r_0_addr[9],
r_2_addr[11]&r_1_addr[3]&r_0_addr[8],
r_2_addr[11]&r_1_addr[3]&r_0_addr[7],
r_2_addr[11]&r_1_addr[3]&r_0_addr[6],
r_2_addr[11]&r_1_addr[3]&r_0_addr[5],
r_2_addr[11]&r_1_addr[3]&r_0_addr[4],
r_2_addr[11]&r_1_addr[3]&r_0_addr[3],
r_2_addr[11]&r_1_addr[3]&r_0_addr[2],
r_2_addr[11]&r_1_addr[3]&r_0_addr[1],
r_2_addr[11]&r_1_addr[3]&r_0_addr[0],
r_2_addr[11]&r_1_addr[2]&r_0_addr[15],
r_2_addr[11]&r_1_addr[2]&r_0_addr[14],
r_2_addr[11]&r_1_addr[2]&r_0_addr[13],
r_2_addr[11]&r_1_addr[2]&r_0_addr[12],
r_2_addr[11]&r_1_addr[2]&r_0_addr[11],
r_2_addr[11]&r_1_addr[2]&r_0_addr[10],
r_2_addr[11]&r_1_addr[2]&r_0_addr[9],
r_2_addr[11]&r_1_addr[2]&r_0_addr[8],
r_2_addr[11]&r_1_addr[2]&r_0_addr[7],
r_2_addr[11]&r_1_addr[2]&r_0_addr[6],
r_2_addr[11]&r_1_addr[2]&r_0_addr[5],
r_2_addr[11]&r_1_addr[2]&r_0_addr[4],
r_2_addr[11]&r_1_addr[2]&r_0_addr[3],
r_2_addr[11]&r_1_addr[2]&r_0_addr[2],
r_2_addr[11]&r_1_addr[2]&r_0_addr[1],
r_2_addr[11]&r_1_addr[2]&r_0_addr[0],
r_2_addr[11]&r_1_addr[1]&r_0_addr[15],
r_2_addr[11]&r_1_addr[1]&r_0_addr[14],
r_2_addr[11]&r_1_addr[1]&r_0_addr[13],
r_2_addr[11]&r_1_addr[1]&r_0_addr[12],
r_2_addr[11]&r_1_addr[1]&r_0_addr[11],
r_2_addr[11]&r_1_addr[1]&r_0_addr[10],
r_2_addr[11]&r_1_addr[1]&r_0_addr[9],
r_2_addr[11]&r_1_addr[1]&r_0_addr[8],
r_2_addr[11]&r_1_addr[1]&r_0_addr[7],
r_2_addr[11]&r_1_addr[1]&r_0_addr[6],
r_2_addr[11]&r_1_addr[1]&r_0_addr[5],
r_2_addr[11]&r_1_addr[1]&r_0_addr[4],
r_2_addr[11]&r_1_addr[1]&r_0_addr[3],
r_2_addr[11]&r_1_addr[1]&r_0_addr[2],
r_2_addr[11]&r_1_addr[1]&r_0_addr[1],
r_2_addr[11]&r_1_addr[1]&r_0_addr[0],
r_2_addr[11]&r_1_addr[0]&r_0_addr[15],
r_2_addr[11]&r_1_addr[0]&r_0_addr[14],
r_2_addr[11]&r_1_addr[0]&r_0_addr[13],
r_2_addr[11]&r_1_addr[0]&r_0_addr[12],
r_2_addr[11]&r_1_addr[0]&r_0_addr[11],
r_2_addr[11]&r_1_addr[0]&r_0_addr[10],
r_2_addr[11]&r_1_addr[0]&r_0_addr[9],
r_2_addr[11]&r_1_addr[0]&r_0_addr[8],
r_2_addr[11]&r_1_addr[0]&r_0_addr[7],
r_2_addr[11]&r_1_addr[0]&r_0_addr[6],
r_2_addr[11]&r_1_addr[0]&r_0_addr[5],
r_2_addr[11]&r_1_addr[0]&r_0_addr[4],
r_2_addr[11]&r_1_addr[0]&r_0_addr[3],
r_2_addr[11]&r_1_addr[0]&r_0_addr[2],
r_2_addr[11]&r_1_addr[0]&r_0_addr[1],
r_2_addr[11]&r_1_addr[0]&r_0_addr[0],
r_2_addr[10]&r_1_addr[15]&r_0_addr[15],
r_2_addr[10]&r_1_addr[15]&r_0_addr[14],
r_2_addr[10]&r_1_addr[15]&r_0_addr[13],
r_2_addr[10]&r_1_addr[15]&r_0_addr[12],
r_2_addr[10]&r_1_addr[15]&r_0_addr[11],
r_2_addr[10]&r_1_addr[15]&r_0_addr[10],
r_2_addr[10]&r_1_addr[15]&r_0_addr[9],
r_2_addr[10]&r_1_addr[15]&r_0_addr[8],
r_2_addr[10]&r_1_addr[15]&r_0_addr[7],
r_2_addr[10]&r_1_addr[15]&r_0_addr[6],
r_2_addr[10]&r_1_addr[15]&r_0_addr[5],
r_2_addr[10]&r_1_addr[15]&r_0_addr[4],
r_2_addr[10]&r_1_addr[15]&r_0_addr[3],
r_2_addr[10]&r_1_addr[15]&r_0_addr[2],
r_2_addr[10]&r_1_addr[15]&r_0_addr[1],
r_2_addr[10]&r_1_addr[15]&r_0_addr[0],
r_2_addr[10]&r_1_addr[14]&r_0_addr[15],
r_2_addr[10]&r_1_addr[14]&r_0_addr[14],
r_2_addr[10]&r_1_addr[14]&r_0_addr[13],
r_2_addr[10]&r_1_addr[14]&r_0_addr[12],
r_2_addr[10]&r_1_addr[14]&r_0_addr[11],
r_2_addr[10]&r_1_addr[14]&r_0_addr[10],
r_2_addr[10]&r_1_addr[14]&r_0_addr[9],
r_2_addr[10]&r_1_addr[14]&r_0_addr[8],
r_2_addr[10]&r_1_addr[14]&r_0_addr[7],
r_2_addr[10]&r_1_addr[14]&r_0_addr[6],
r_2_addr[10]&r_1_addr[14]&r_0_addr[5],
r_2_addr[10]&r_1_addr[14]&r_0_addr[4],
r_2_addr[10]&r_1_addr[14]&r_0_addr[3],
r_2_addr[10]&r_1_addr[14]&r_0_addr[2],
r_2_addr[10]&r_1_addr[14]&r_0_addr[1],
r_2_addr[10]&r_1_addr[14]&r_0_addr[0],
r_2_addr[10]&r_1_addr[13]&r_0_addr[15],
r_2_addr[10]&r_1_addr[13]&r_0_addr[14],
r_2_addr[10]&r_1_addr[13]&r_0_addr[13],
r_2_addr[10]&r_1_addr[13]&r_0_addr[12],
r_2_addr[10]&r_1_addr[13]&r_0_addr[11],
r_2_addr[10]&r_1_addr[13]&r_0_addr[10],
r_2_addr[10]&r_1_addr[13]&r_0_addr[9],
r_2_addr[10]&r_1_addr[13]&r_0_addr[8],
r_2_addr[10]&r_1_addr[13]&r_0_addr[7],
r_2_addr[10]&r_1_addr[13]&r_0_addr[6],
r_2_addr[10]&r_1_addr[13]&r_0_addr[5],
r_2_addr[10]&r_1_addr[13]&r_0_addr[4],
r_2_addr[10]&r_1_addr[13]&r_0_addr[3],
r_2_addr[10]&r_1_addr[13]&r_0_addr[2],
r_2_addr[10]&r_1_addr[13]&r_0_addr[1],
r_2_addr[10]&r_1_addr[13]&r_0_addr[0],
r_2_addr[10]&r_1_addr[12]&r_0_addr[15],
r_2_addr[10]&r_1_addr[12]&r_0_addr[14],
r_2_addr[10]&r_1_addr[12]&r_0_addr[13],
r_2_addr[10]&r_1_addr[12]&r_0_addr[12],
r_2_addr[10]&r_1_addr[12]&r_0_addr[11],
r_2_addr[10]&r_1_addr[12]&r_0_addr[10],
r_2_addr[10]&r_1_addr[12]&r_0_addr[9],
r_2_addr[10]&r_1_addr[12]&r_0_addr[8],
r_2_addr[10]&r_1_addr[12]&r_0_addr[7],
r_2_addr[10]&r_1_addr[12]&r_0_addr[6],
r_2_addr[10]&r_1_addr[12]&r_0_addr[5],
r_2_addr[10]&r_1_addr[12]&r_0_addr[4],
r_2_addr[10]&r_1_addr[12]&r_0_addr[3],
r_2_addr[10]&r_1_addr[12]&r_0_addr[2],
r_2_addr[10]&r_1_addr[12]&r_0_addr[1],
r_2_addr[10]&r_1_addr[12]&r_0_addr[0],
r_2_addr[10]&r_1_addr[11]&r_0_addr[15],
r_2_addr[10]&r_1_addr[11]&r_0_addr[14],
r_2_addr[10]&r_1_addr[11]&r_0_addr[13],
r_2_addr[10]&r_1_addr[11]&r_0_addr[12],
r_2_addr[10]&r_1_addr[11]&r_0_addr[11],
r_2_addr[10]&r_1_addr[11]&r_0_addr[10],
r_2_addr[10]&r_1_addr[11]&r_0_addr[9],
r_2_addr[10]&r_1_addr[11]&r_0_addr[8],
r_2_addr[10]&r_1_addr[11]&r_0_addr[7],
r_2_addr[10]&r_1_addr[11]&r_0_addr[6],
r_2_addr[10]&r_1_addr[11]&r_0_addr[5],
r_2_addr[10]&r_1_addr[11]&r_0_addr[4],
r_2_addr[10]&r_1_addr[11]&r_0_addr[3],
r_2_addr[10]&r_1_addr[11]&r_0_addr[2],
r_2_addr[10]&r_1_addr[11]&r_0_addr[1],
r_2_addr[10]&r_1_addr[11]&r_0_addr[0],
r_2_addr[10]&r_1_addr[10]&r_0_addr[15],
r_2_addr[10]&r_1_addr[10]&r_0_addr[14],
r_2_addr[10]&r_1_addr[10]&r_0_addr[13],
r_2_addr[10]&r_1_addr[10]&r_0_addr[12],
r_2_addr[10]&r_1_addr[10]&r_0_addr[11],
r_2_addr[10]&r_1_addr[10]&r_0_addr[10],
r_2_addr[10]&r_1_addr[10]&r_0_addr[9],
r_2_addr[10]&r_1_addr[10]&r_0_addr[8],
r_2_addr[10]&r_1_addr[10]&r_0_addr[7],
r_2_addr[10]&r_1_addr[10]&r_0_addr[6],
r_2_addr[10]&r_1_addr[10]&r_0_addr[5],
r_2_addr[10]&r_1_addr[10]&r_0_addr[4],
r_2_addr[10]&r_1_addr[10]&r_0_addr[3],
r_2_addr[10]&r_1_addr[10]&r_0_addr[2],
r_2_addr[10]&r_1_addr[10]&r_0_addr[1],
r_2_addr[10]&r_1_addr[10]&r_0_addr[0],
r_2_addr[10]&r_1_addr[9]&r_0_addr[15],
r_2_addr[10]&r_1_addr[9]&r_0_addr[14],
r_2_addr[10]&r_1_addr[9]&r_0_addr[13],
r_2_addr[10]&r_1_addr[9]&r_0_addr[12],
r_2_addr[10]&r_1_addr[9]&r_0_addr[11],
r_2_addr[10]&r_1_addr[9]&r_0_addr[10],
r_2_addr[10]&r_1_addr[9]&r_0_addr[9],
r_2_addr[10]&r_1_addr[9]&r_0_addr[8],
r_2_addr[10]&r_1_addr[9]&r_0_addr[7],
r_2_addr[10]&r_1_addr[9]&r_0_addr[6],
r_2_addr[10]&r_1_addr[9]&r_0_addr[5],
r_2_addr[10]&r_1_addr[9]&r_0_addr[4],
r_2_addr[10]&r_1_addr[9]&r_0_addr[3],
r_2_addr[10]&r_1_addr[9]&r_0_addr[2],
r_2_addr[10]&r_1_addr[9]&r_0_addr[1],
r_2_addr[10]&r_1_addr[9]&r_0_addr[0],
r_2_addr[10]&r_1_addr[8]&r_0_addr[15],
r_2_addr[10]&r_1_addr[8]&r_0_addr[14],
r_2_addr[10]&r_1_addr[8]&r_0_addr[13],
r_2_addr[10]&r_1_addr[8]&r_0_addr[12],
r_2_addr[10]&r_1_addr[8]&r_0_addr[11],
r_2_addr[10]&r_1_addr[8]&r_0_addr[10],
r_2_addr[10]&r_1_addr[8]&r_0_addr[9],
r_2_addr[10]&r_1_addr[8]&r_0_addr[8],
r_2_addr[10]&r_1_addr[8]&r_0_addr[7],
r_2_addr[10]&r_1_addr[8]&r_0_addr[6],
r_2_addr[10]&r_1_addr[8]&r_0_addr[5],
r_2_addr[10]&r_1_addr[8]&r_0_addr[4],
r_2_addr[10]&r_1_addr[8]&r_0_addr[3],
r_2_addr[10]&r_1_addr[8]&r_0_addr[2],
r_2_addr[10]&r_1_addr[8]&r_0_addr[1],
r_2_addr[10]&r_1_addr[8]&r_0_addr[0],
r_2_addr[10]&r_1_addr[7]&r_0_addr[15],
r_2_addr[10]&r_1_addr[7]&r_0_addr[14],
r_2_addr[10]&r_1_addr[7]&r_0_addr[13],
r_2_addr[10]&r_1_addr[7]&r_0_addr[12],
r_2_addr[10]&r_1_addr[7]&r_0_addr[11],
r_2_addr[10]&r_1_addr[7]&r_0_addr[10],
r_2_addr[10]&r_1_addr[7]&r_0_addr[9],
r_2_addr[10]&r_1_addr[7]&r_0_addr[8],
r_2_addr[10]&r_1_addr[7]&r_0_addr[7],
r_2_addr[10]&r_1_addr[7]&r_0_addr[6],
r_2_addr[10]&r_1_addr[7]&r_0_addr[5],
r_2_addr[10]&r_1_addr[7]&r_0_addr[4],
r_2_addr[10]&r_1_addr[7]&r_0_addr[3],
r_2_addr[10]&r_1_addr[7]&r_0_addr[2],
r_2_addr[10]&r_1_addr[7]&r_0_addr[1],
r_2_addr[10]&r_1_addr[7]&r_0_addr[0],
r_2_addr[10]&r_1_addr[6]&r_0_addr[15],
r_2_addr[10]&r_1_addr[6]&r_0_addr[14],
r_2_addr[10]&r_1_addr[6]&r_0_addr[13],
r_2_addr[10]&r_1_addr[6]&r_0_addr[12],
r_2_addr[10]&r_1_addr[6]&r_0_addr[11],
r_2_addr[10]&r_1_addr[6]&r_0_addr[10],
r_2_addr[10]&r_1_addr[6]&r_0_addr[9],
r_2_addr[10]&r_1_addr[6]&r_0_addr[8],
r_2_addr[10]&r_1_addr[6]&r_0_addr[7],
r_2_addr[10]&r_1_addr[6]&r_0_addr[6],
r_2_addr[10]&r_1_addr[6]&r_0_addr[5],
r_2_addr[10]&r_1_addr[6]&r_0_addr[4],
r_2_addr[10]&r_1_addr[6]&r_0_addr[3],
r_2_addr[10]&r_1_addr[6]&r_0_addr[2],
r_2_addr[10]&r_1_addr[6]&r_0_addr[1],
r_2_addr[10]&r_1_addr[6]&r_0_addr[0],
r_2_addr[10]&r_1_addr[5]&r_0_addr[15],
r_2_addr[10]&r_1_addr[5]&r_0_addr[14],
r_2_addr[10]&r_1_addr[5]&r_0_addr[13],
r_2_addr[10]&r_1_addr[5]&r_0_addr[12],
r_2_addr[10]&r_1_addr[5]&r_0_addr[11],
r_2_addr[10]&r_1_addr[5]&r_0_addr[10],
r_2_addr[10]&r_1_addr[5]&r_0_addr[9],
r_2_addr[10]&r_1_addr[5]&r_0_addr[8],
r_2_addr[10]&r_1_addr[5]&r_0_addr[7],
r_2_addr[10]&r_1_addr[5]&r_0_addr[6],
r_2_addr[10]&r_1_addr[5]&r_0_addr[5],
r_2_addr[10]&r_1_addr[5]&r_0_addr[4],
r_2_addr[10]&r_1_addr[5]&r_0_addr[3],
r_2_addr[10]&r_1_addr[5]&r_0_addr[2],
r_2_addr[10]&r_1_addr[5]&r_0_addr[1],
r_2_addr[10]&r_1_addr[5]&r_0_addr[0],
r_2_addr[10]&r_1_addr[4]&r_0_addr[15],
r_2_addr[10]&r_1_addr[4]&r_0_addr[14],
r_2_addr[10]&r_1_addr[4]&r_0_addr[13],
r_2_addr[10]&r_1_addr[4]&r_0_addr[12],
r_2_addr[10]&r_1_addr[4]&r_0_addr[11],
r_2_addr[10]&r_1_addr[4]&r_0_addr[10],
r_2_addr[10]&r_1_addr[4]&r_0_addr[9],
r_2_addr[10]&r_1_addr[4]&r_0_addr[8],
r_2_addr[10]&r_1_addr[4]&r_0_addr[7],
r_2_addr[10]&r_1_addr[4]&r_0_addr[6],
r_2_addr[10]&r_1_addr[4]&r_0_addr[5],
r_2_addr[10]&r_1_addr[4]&r_0_addr[4],
r_2_addr[10]&r_1_addr[4]&r_0_addr[3],
r_2_addr[10]&r_1_addr[4]&r_0_addr[2],
r_2_addr[10]&r_1_addr[4]&r_0_addr[1],
r_2_addr[10]&r_1_addr[4]&r_0_addr[0],
r_2_addr[10]&r_1_addr[3]&r_0_addr[15],
r_2_addr[10]&r_1_addr[3]&r_0_addr[14],
r_2_addr[10]&r_1_addr[3]&r_0_addr[13],
r_2_addr[10]&r_1_addr[3]&r_0_addr[12],
r_2_addr[10]&r_1_addr[3]&r_0_addr[11],
r_2_addr[10]&r_1_addr[3]&r_0_addr[10],
r_2_addr[10]&r_1_addr[3]&r_0_addr[9],
r_2_addr[10]&r_1_addr[3]&r_0_addr[8],
r_2_addr[10]&r_1_addr[3]&r_0_addr[7],
r_2_addr[10]&r_1_addr[3]&r_0_addr[6],
r_2_addr[10]&r_1_addr[3]&r_0_addr[5],
r_2_addr[10]&r_1_addr[3]&r_0_addr[4],
r_2_addr[10]&r_1_addr[3]&r_0_addr[3],
r_2_addr[10]&r_1_addr[3]&r_0_addr[2],
r_2_addr[10]&r_1_addr[3]&r_0_addr[1],
r_2_addr[10]&r_1_addr[3]&r_0_addr[0],
r_2_addr[10]&r_1_addr[2]&r_0_addr[15],
r_2_addr[10]&r_1_addr[2]&r_0_addr[14],
r_2_addr[10]&r_1_addr[2]&r_0_addr[13],
r_2_addr[10]&r_1_addr[2]&r_0_addr[12],
r_2_addr[10]&r_1_addr[2]&r_0_addr[11],
r_2_addr[10]&r_1_addr[2]&r_0_addr[10],
r_2_addr[10]&r_1_addr[2]&r_0_addr[9],
r_2_addr[10]&r_1_addr[2]&r_0_addr[8],
r_2_addr[10]&r_1_addr[2]&r_0_addr[7],
r_2_addr[10]&r_1_addr[2]&r_0_addr[6],
r_2_addr[10]&r_1_addr[2]&r_0_addr[5],
r_2_addr[10]&r_1_addr[2]&r_0_addr[4],
r_2_addr[10]&r_1_addr[2]&r_0_addr[3],
r_2_addr[10]&r_1_addr[2]&r_0_addr[2],
r_2_addr[10]&r_1_addr[2]&r_0_addr[1],
r_2_addr[10]&r_1_addr[2]&r_0_addr[0],
r_2_addr[10]&r_1_addr[1]&r_0_addr[15],
r_2_addr[10]&r_1_addr[1]&r_0_addr[14],
r_2_addr[10]&r_1_addr[1]&r_0_addr[13],
r_2_addr[10]&r_1_addr[1]&r_0_addr[12],
r_2_addr[10]&r_1_addr[1]&r_0_addr[11],
r_2_addr[10]&r_1_addr[1]&r_0_addr[10],
r_2_addr[10]&r_1_addr[1]&r_0_addr[9],
r_2_addr[10]&r_1_addr[1]&r_0_addr[8],
r_2_addr[10]&r_1_addr[1]&r_0_addr[7],
r_2_addr[10]&r_1_addr[1]&r_0_addr[6],
r_2_addr[10]&r_1_addr[1]&r_0_addr[5],
r_2_addr[10]&r_1_addr[1]&r_0_addr[4],
r_2_addr[10]&r_1_addr[1]&r_0_addr[3],
r_2_addr[10]&r_1_addr[1]&r_0_addr[2],
r_2_addr[10]&r_1_addr[1]&r_0_addr[1],
r_2_addr[10]&r_1_addr[1]&r_0_addr[0],
r_2_addr[10]&r_1_addr[0]&r_0_addr[15],
r_2_addr[10]&r_1_addr[0]&r_0_addr[14],
r_2_addr[10]&r_1_addr[0]&r_0_addr[13],
r_2_addr[10]&r_1_addr[0]&r_0_addr[12],
r_2_addr[10]&r_1_addr[0]&r_0_addr[11],
r_2_addr[10]&r_1_addr[0]&r_0_addr[10],
r_2_addr[10]&r_1_addr[0]&r_0_addr[9],
r_2_addr[10]&r_1_addr[0]&r_0_addr[8],
r_2_addr[10]&r_1_addr[0]&r_0_addr[7],
r_2_addr[10]&r_1_addr[0]&r_0_addr[6],
r_2_addr[10]&r_1_addr[0]&r_0_addr[5],
r_2_addr[10]&r_1_addr[0]&r_0_addr[4],
r_2_addr[10]&r_1_addr[0]&r_0_addr[3],
r_2_addr[10]&r_1_addr[0]&r_0_addr[2],
r_2_addr[10]&r_1_addr[0]&r_0_addr[1],
r_2_addr[10]&r_1_addr[0]&r_0_addr[0],
r_2_addr[9]&r_1_addr[15]&r_0_addr[15],
r_2_addr[9]&r_1_addr[15]&r_0_addr[14],
r_2_addr[9]&r_1_addr[15]&r_0_addr[13],
r_2_addr[9]&r_1_addr[15]&r_0_addr[12],
r_2_addr[9]&r_1_addr[15]&r_0_addr[11],
r_2_addr[9]&r_1_addr[15]&r_0_addr[10],
r_2_addr[9]&r_1_addr[15]&r_0_addr[9],
r_2_addr[9]&r_1_addr[15]&r_0_addr[8],
r_2_addr[9]&r_1_addr[15]&r_0_addr[7],
r_2_addr[9]&r_1_addr[15]&r_0_addr[6],
r_2_addr[9]&r_1_addr[15]&r_0_addr[5],
r_2_addr[9]&r_1_addr[15]&r_0_addr[4],
r_2_addr[9]&r_1_addr[15]&r_0_addr[3],
r_2_addr[9]&r_1_addr[15]&r_0_addr[2],
r_2_addr[9]&r_1_addr[15]&r_0_addr[1],
r_2_addr[9]&r_1_addr[15]&r_0_addr[0],
r_2_addr[9]&r_1_addr[14]&r_0_addr[15],
r_2_addr[9]&r_1_addr[14]&r_0_addr[14],
r_2_addr[9]&r_1_addr[14]&r_0_addr[13],
r_2_addr[9]&r_1_addr[14]&r_0_addr[12],
r_2_addr[9]&r_1_addr[14]&r_0_addr[11],
r_2_addr[9]&r_1_addr[14]&r_0_addr[10],
r_2_addr[9]&r_1_addr[14]&r_0_addr[9],
r_2_addr[9]&r_1_addr[14]&r_0_addr[8],
r_2_addr[9]&r_1_addr[14]&r_0_addr[7],
r_2_addr[9]&r_1_addr[14]&r_0_addr[6],
r_2_addr[9]&r_1_addr[14]&r_0_addr[5],
r_2_addr[9]&r_1_addr[14]&r_0_addr[4],
r_2_addr[9]&r_1_addr[14]&r_0_addr[3],
r_2_addr[9]&r_1_addr[14]&r_0_addr[2],
r_2_addr[9]&r_1_addr[14]&r_0_addr[1],
r_2_addr[9]&r_1_addr[14]&r_0_addr[0],
r_2_addr[9]&r_1_addr[13]&r_0_addr[15],
r_2_addr[9]&r_1_addr[13]&r_0_addr[14],
r_2_addr[9]&r_1_addr[13]&r_0_addr[13],
r_2_addr[9]&r_1_addr[13]&r_0_addr[12],
r_2_addr[9]&r_1_addr[13]&r_0_addr[11],
r_2_addr[9]&r_1_addr[13]&r_0_addr[10],
r_2_addr[9]&r_1_addr[13]&r_0_addr[9],
r_2_addr[9]&r_1_addr[13]&r_0_addr[8],
r_2_addr[9]&r_1_addr[13]&r_0_addr[7],
r_2_addr[9]&r_1_addr[13]&r_0_addr[6],
r_2_addr[9]&r_1_addr[13]&r_0_addr[5],
r_2_addr[9]&r_1_addr[13]&r_0_addr[4],
r_2_addr[9]&r_1_addr[13]&r_0_addr[3],
r_2_addr[9]&r_1_addr[13]&r_0_addr[2],
r_2_addr[9]&r_1_addr[13]&r_0_addr[1],
r_2_addr[9]&r_1_addr[13]&r_0_addr[0],
r_2_addr[9]&r_1_addr[12]&r_0_addr[15],
r_2_addr[9]&r_1_addr[12]&r_0_addr[14],
r_2_addr[9]&r_1_addr[12]&r_0_addr[13],
r_2_addr[9]&r_1_addr[12]&r_0_addr[12],
r_2_addr[9]&r_1_addr[12]&r_0_addr[11],
r_2_addr[9]&r_1_addr[12]&r_0_addr[10],
r_2_addr[9]&r_1_addr[12]&r_0_addr[9],
r_2_addr[9]&r_1_addr[12]&r_0_addr[8],
r_2_addr[9]&r_1_addr[12]&r_0_addr[7],
r_2_addr[9]&r_1_addr[12]&r_0_addr[6],
r_2_addr[9]&r_1_addr[12]&r_0_addr[5],
r_2_addr[9]&r_1_addr[12]&r_0_addr[4],
r_2_addr[9]&r_1_addr[12]&r_0_addr[3],
r_2_addr[9]&r_1_addr[12]&r_0_addr[2],
r_2_addr[9]&r_1_addr[12]&r_0_addr[1],
r_2_addr[9]&r_1_addr[12]&r_0_addr[0],
r_2_addr[9]&r_1_addr[11]&r_0_addr[15],
r_2_addr[9]&r_1_addr[11]&r_0_addr[14],
r_2_addr[9]&r_1_addr[11]&r_0_addr[13],
r_2_addr[9]&r_1_addr[11]&r_0_addr[12],
r_2_addr[9]&r_1_addr[11]&r_0_addr[11],
r_2_addr[9]&r_1_addr[11]&r_0_addr[10],
r_2_addr[9]&r_1_addr[11]&r_0_addr[9],
r_2_addr[9]&r_1_addr[11]&r_0_addr[8],
r_2_addr[9]&r_1_addr[11]&r_0_addr[7],
r_2_addr[9]&r_1_addr[11]&r_0_addr[6],
r_2_addr[9]&r_1_addr[11]&r_0_addr[5],
r_2_addr[9]&r_1_addr[11]&r_0_addr[4],
r_2_addr[9]&r_1_addr[11]&r_0_addr[3],
r_2_addr[9]&r_1_addr[11]&r_0_addr[2],
r_2_addr[9]&r_1_addr[11]&r_0_addr[1],
r_2_addr[9]&r_1_addr[11]&r_0_addr[0],
r_2_addr[9]&r_1_addr[10]&r_0_addr[15],
r_2_addr[9]&r_1_addr[10]&r_0_addr[14],
r_2_addr[9]&r_1_addr[10]&r_0_addr[13],
r_2_addr[9]&r_1_addr[10]&r_0_addr[12],
r_2_addr[9]&r_1_addr[10]&r_0_addr[11],
r_2_addr[9]&r_1_addr[10]&r_0_addr[10],
r_2_addr[9]&r_1_addr[10]&r_0_addr[9],
r_2_addr[9]&r_1_addr[10]&r_0_addr[8],
r_2_addr[9]&r_1_addr[10]&r_0_addr[7],
r_2_addr[9]&r_1_addr[10]&r_0_addr[6],
r_2_addr[9]&r_1_addr[10]&r_0_addr[5],
r_2_addr[9]&r_1_addr[10]&r_0_addr[4],
r_2_addr[9]&r_1_addr[10]&r_0_addr[3],
r_2_addr[9]&r_1_addr[10]&r_0_addr[2],
r_2_addr[9]&r_1_addr[10]&r_0_addr[1],
r_2_addr[9]&r_1_addr[10]&r_0_addr[0],
r_2_addr[9]&r_1_addr[9]&r_0_addr[15],
r_2_addr[9]&r_1_addr[9]&r_0_addr[14],
r_2_addr[9]&r_1_addr[9]&r_0_addr[13],
r_2_addr[9]&r_1_addr[9]&r_0_addr[12],
r_2_addr[9]&r_1_addr[9]&r_0_addr[11],
r_2_addr[9]&r_1_addr[9]&r_0_addr[10],
r_2_addr[9]&r_1_addr[9]&r_0_addr[9],
r_2_addr[9]&r_1_addr[9]&r_0_addr[8],
r_2_addr[9]&r_1_addr[9]&r_0_addr[7],
r_2_addr[9]&r_1_addr[9]&r_0_addr[6],
r_2_addr[9]&r_1_addr[9]&r_0_addr[5],
r_2_addr[9]&r_1_addr[9]&r_0_addr[4],
r_2_addr[9]&r_1_addr[9]&r_0_addr[3],
r_2_addr[9]&r_1_addr[9]&r_0_addr[2],
r_2_addr[9]&r_1_addr[9]&r_0_addr[1],
r_2_addr[9]&r_1_addr[9]&r_0_addr[0],
r_2_addr[9]&r_1_addr[8]&r_0_addr[15],
r_2_addr[9]&r_1_addr[8]&r_0_addr[14],
r_2_addr[9]&r_1_addr[8]&r_0_addr[13],
r_2_addr[9]&r_1_addr[8]&r_0_addr[12],
r_2_addr[9]&r_1_addr[8]&r_0_addr[11],
r_2_addr[9]&r_1_addr[8]&r_0_addr[10],
r_2_addr[9]&r_1_addr[8]&r_0_addr[9],
r_2_addr[9]&r_1_addr[8]&r_0_addr[8],
r_2_addr[9]&r_1_addr[8]&r_0_addr[7],
r_2_addr[9]&r_1_addr[8]&r_0_addr[6],
r_2_addr[9]&r_1_addr[8]&r_0_addr[5],
r_2_addr[9]&r_1_addr[8]&r_0_addr[4],
r_2_addr[9]&r_1_addr[8]&r_0_addr[3],
r_2_addr[9]&r_1_addr[8]&r_0_addr[2],
r_2_addr[9]&r_1_addr[8]&r_0_addr[1],
r_2_addr[9]&r_1_addr[8]&r_0_addr[0],
r_2_addr[9]&r_1_addr[7]&r_0_addr[15],
r_2_addr[9]&r_1_addr[7]&r_0_addr[14],
r_2_addr[9]&r_1_addr[7]&r_0_addr[13],
r_2_addr[9]&r_1_addr[7]&r_0_addr[12],
r_2_addr[9]&r_1_addr[7]&r_0_addr[11],
r_2_addr[9]&r_1_addr[7]&r_0_addr[10],
r_2_addr[9]&r_1_addr[7]&r_0_addr[9],
r_2_addr[9]&r_1_addr[7]&r_0_addr[8],
r_2_addr[9]&r_1_addr[7]&r_0_addr[7],
r_2_addr[9]&r_1_addr[7]&r_0_addr[6],
r_2_addr[9]&r_1_addr[7]&r_0_addr[5],
r_2_addr[9]&r_1_addr[7]&r_0_addr[4],
r_2_addr[9]&r_1_addr[7]&r_0_addr[3],
r_2_addr[9]&r_1_addr[7]&r_0_addr[2],
r_2_addr[9]&r_1_addr[7]&r_0_addr[1],
r_2_addr[9]&r_1_addr[7]&r_0_addr[0],
r_2_addr[9]&r_1_addr[6]&r_0_addr[15],
r_2_addr[9]&r_1_addr[6]&r_0_addr[14],
r_2_addr[9]&r_1_addr[6]&r_0_addr[13],
r_2_addr[9]&r_1_addr[6]&r_0_addr[12],
r_2_addr[9]&r_1_addr[6]&r_0_addr[11],
r_2_addr[9]&r_1_addr[6]&r_0_addr[10],
r_2_addr[9]&r_1_addr[6]&r_0_addr[9],
r_2_addr[9]&r_1_addr[6]&r_0_addr[8],
r_2_addr[9]&r_1_addr[6]&r_0_addr[7],
r_2_addr[9]&r_1_addr[6]&r_0_addr[6],
r_2_addr[9]&r_1_addr[6]&r_0_addr[5],
r_2_addr[9]&r_1_addr[6]&r_0_addr[4],
r_2_addr[9]&r_1_addr[6]&r_0_addr[3],
r_2_addr[9]&r_1_addr[6]&r_0_addr[2],
r_2_addr[9]&r_1_addr[6]&r_0_addr[1],
r_2_addr[9]&r_1_addr[6]&r_0_addr[0],
r_2_addr[9]&r_1_addr[5]&r_0_addr[15],
r_2_addr[9]&r_1_addr[5]&r_0_addr[14],
r_2_addr[9]&r_1_addr[5]&r_0_addr[13],
r_2_addr[9]&r_1_addr[5]&r_0_addr[12],
r_2_addr[9]&r_1_addr[5]&r_0_addr[11],
r_2_addr[9]&r_1_addr[5]&r_0_addr[10],
r_2_addr[9]&r_1_addr[5]&r_0_addr[9],
r_2_addr[9]&r_1_addr[5]&r_0_addr[8],
r_2_addr[9]&r_1_addr[5]&r_0_addr[7],
r_2_addr[9]&r_1_addr[5]&r_0_addr[6],
r_2_addr[9]&r_1_addr[5]&r_0_addr[5],
r_2_addr[9]&r_1_addr[5]&r_0_addr[4],
r_2_addr[9]&r_1_addr[5]&r_0_addr[3],
r_2_addr[9]&r_1_addr[5]&r_0_addr[2],
r_2_addr[9]&r_1_addr[5]&r_0_addr[1],
r_2_addr[9]&r_1_addr[5]&r_0_addr[0],
r_2_addr[9]&r_1_addr[4]&r_0_addr[15],
r_2_addr[9]&r_1_addr[4]&r_0_addr[14],
r_2_addr[9]&r_1_addr[4]&r_0_addr[13],
r_2_addr[9]&r_1_addr[4]&r_0_addr[12],
r_2_addr[9]&r_1_addr[4]&r_0_addr[11],
r_2_addr[9]&r_1_addr[4]&r_0_addr[10],
r_2_addr[9]&r_1_addr[4]&r_0_addr[9],
r_2_addr[9]&r_1_addr[4]&r_0_addr[8],
r_2_addr[9]&r_1_addr[4]&r_0_addr[7],
r_2_addr[9]&r_1_addr[4]&r_0_addr[6],
r_2_addr[9]&r_1_addr[4]&r_0_addr[5],
r_2_addr[9]&r_1_addr[4]&r_0_addr[4],
r_2_addr[9]&r_1_addr[4]&r_0_addr[3],
r_2_addr[9]&r_1_addr[4]&r_0_addr[2],
r_2_addr[9]&r_1_addr[4]&r_0_addr[1],
r_2_addr[9]&r_1_addr[4]&r_0_addr[0],
r_2_addr[9]&r_1_addr[3]&r_0_addr[15],
r_2_addr[9]&r_1_addr[3]&r_0_addr[14],
r_2_addr[9]&r_1_addr[3]&r_0_addr[13],
r_2_addr[9]&r_1_addr[3]&r_0_addr[12],
r_2_addr[9]&r_1_addr[3]&r_0_addr[11],
r_2_addr[9]&r_1_addr[3]&r_0_addr[10],
r_2_addr[9]&r_1_addr[3]&r_0_addr[9],
r_2_addr[9]&r_1_addr[3]&r_0_addr[8],
r_2_addr[9]&r_1_addr[3]&r_0_addr[7],
r_2_addr[9]&r_1_addr[3]&r_0_addr[6],
r_2_addr[9]&r_1_addr[3]&r_0_addr[5],
r_2_addr[9]&r_1_addr[3]&r_0_addr[4],
r_2_addr[9]&r_1_addr[3]&r_0_addr[3],
r_2_addr[9]&r_1_addr[3]&r_0_addr[2],
r_2_addr[9]&r_1_addr[3]&r_0_addr[1],
r_2_addr[9]&r_1_addr[3]&r_0_addr[0],
r_2_addr[9]&r_1_addr[2]&r_0_addr[15],
r_2_addr[9]&r_1_addr[2]&r_0_addr[14],
r_2_addr[9]&r_1_addr[2]&r_0_addr[13],
r_2_addr[9]&r_1_addr[2]&r_0_addr[12],
r_2_addr[9]&r_1_addr[2]&r_0_addr[11],
r_2_addr[9]&r_1_addr[2]&r_0_addr[10],
r_2_addr[9]&r_1_addr[2]&r_0_addr[9],
r_2_addr[9]&r_1_addr[2]&r_0_addr[8],
r_2_addr[9]&r_1_addr[2]&r_0_addr[7],
r_2_addr[9]&r_1_addr[2]&r_0_addr[6],
r_2_addr[9]&r_1_addr[2]&r_0_addr[5],
r_2_addr[9]&r_1_addr[2]&r_0_addr[4],
r_2_addr[9]&r_1_addr[2]&r_0_addr[3],
r_2_addr[9]&r_1_addr[2]&r_0_addr[2],
r_2_addr[9]&r_1_addr[2]&r_0_addr[1],
r_2_addr[9]&r_1_addr[2]&r_0_addr[0],
r_2_addr[9]&r_1_addr[1]&r_0_addr[15],
r_2_addr[9]&r_1_addr[1]&r_0_addr[14],
r_2_addr[9]&r_1_addr[1]&r_0_addr[13],
r_2_addr[9]&r_1_addr[1]&r_0_addr[12],
r_2_addr[9]&r_1_addr[1]&r_0_addr[11],
r_2_addr[9]&r_1_addr[1]&r_0_addr[10],
r_2_addr[9]&r_1_addr[1]&r_0_addr[9],
r_2_addr[9]&r_1_addr[1]&r_0_addr[8],
r_2_addr[9]&r_1_addr[1]&r_0_addr[7],
r_2_addr[9]&r_1_addr[1]&r_0_addr[6],
r_2_addr[9]&r_1_addr[1]&r_0_addr[5],
r_2_addr[9]&r_1_addr[1]&r_0_addr[4],
r_2_addr[9]&r_1_addr[1]&r_0_addr[3],
r_2_addr[9]&r_1_addr[1]&r_0_addr[2],
r_2_addr[9]&r_1_addr[1]&r_0_addr[1],
r_2_addr[9]&r_1_addr[1]&r_0_addr[0],
r_2_addr[9]&r_1_addr[0]&r_0_addr[15],
r_2_addr[9]&r_1_addr[0]&r_0_addr[14],
r_2_addr[9]&r_1_addr[0]&r_0_addr[13],
r_2_addr[9]&r_1_addr[0]&r_0_addr[12],
r_2_addr[9]&r_1_addr[0]&r_0_addr[11],
r_2_addr[9]&r_1_addr[0]&r_0_addr[10],
r_2_addr[9]&r_1_addr[0]&r_0_addr[9],
r_2_addr[9]&r_1_addr[0]&r_0_addr[8],
r_2_addr[9]&r_1_addr[0]&r_0_addr[7],
r_2_addr[9]&r_1_addr[0]&r_0_addr[6],
r_2_addr[9]&r_1_addr[0]&r_0_addr[5],
r_2_addr[9]&r_1_addr[0]&r_0_addr[4],
r_2_addr[9]&r_1_addr[0]&r_0_addr[3],
r_2_addr[9]&r_1_addr[0]&r_0_addr[2],
r_2_addr[9]&r_1_addr[0]&r_0_addr[1],
r_2_addr[9]&r_1_addr[0]&r_0_addr[0],
r_2_addr[8]&r_1_addr[15]&r_0_addr[15],
r_2_addr[8]&r_1_addr[15]&r_0_addr[14],
r_2_addr[8]&r_1_addr[15]&r_0_addr[13],
r_2_addr[8]&r_1_addr[15]&r_0_addr[12],
r_2_addr[8]&r_1_addr[15]&r_0_addr[11],
r_2_addr[8]&r_1_addr[15]&r_0_addr[10],
r_2_addr[8]&r_1_addr[15]&r_0_addr[9],
r_2_addr[8]&r_1_addr[15]&r_0_addr[8],
r_2_addr[8]&r_1_addr[15]&r_0_addr[7],
r_2_addr[8]&r_1_addr[15]&r_0_addr[6],
r_2_addr[8]&r_1_addr[15]&r_0_addr[5],
r_2_addr[8]&r_1_addr[15]&r_0_addr[4],
r_2_addr[8]&r_1_addr[15]&r_0_addr[3],
r_2_addr[8]&r_1_addr[15]&r_0_addr[2],
r_2_addr[8]&r_1_addr[15]&r_0_addr[1],
r_2_addr[8]&r_1_addr[15]&r_0_addr[0],
r_2_addr[8]&r_1_addr[14]&r_0_addr[15],
r_2_addr[8]&r_1_addr[14]&r_0_addr[14],
r_2_addr[8]&r_1_addr[14]&r_0_addr[13],
r_2_addr[8]&r_1_addr[14]&r_0_addr[12],
r_2_addr[8]&r_1_addr[14]&r_0_addr[11],
r_2_addr[8]&r_1_addr[14]&r_0_addr[10],
r_2_addr[8]&r_1_addr[14]&r_0_addr[9],
r_2_addr[8]&r_1_addr[14]&r_0_addr[8],
r_2_addr[8]&r_1_addr[14]&r_0_addr[7],
r_2_addr[8]&r_1_addr[14]&r_0_addr[6],
r_2_addr[8]&r_1_addr[14]&r_0_addr[5],
r_2_addr[8]&r_1_addr[14]&r_0_addr[4],
r_2_addr[8]&r_1_addr[14]&r_0_addr[3],
r_2_addr[8]&r_1_addr[14]&r_0_addr[2],
r_2_addr[8]&r_1_addr[14]&r_0_addr[1],
r_2_addr[8]&r_1_addr[14]&r_0_addr[0],
r_2_addr[8]&r_1_addr[13]&r_0_addr[15],
r_2_addr[8]&r_1_addr[13]&r_0_addr[14],
r_2_addr[8]&r_1_addr[13]&r_0_addr[13],
r_2_addr[8]&r_1_addr[13]&r_0_addr[12],
r_2_addr[8]&r_1_addr[13]&r_0_addr[11],
r_2_addr[8]&r_1_addr[13]&r_0_addr[10],
r_2_addr[8]&r_1_addr[13]&r_0_addr[9],
r_2_addr[8]&r_1_addr[13]&r_0_addr[8],
r_2_addr[8]&r_1_addr[13]&r_0_addr[7],
r_2_addr[8]&r_1_addr[13]&r_0_addr[6],
r_2_addr[8]&r_1_addr[13]&r_0_addr[5],
r_2_addr[8]&r_1_addr[13]&r_0_addr[4],
r_2_addr[8]&r_1_addr[13]&r_0_addr[3],
r_2_addr[8]&r_1_addr[13]&r_0_addr[2],
r_2_addr[8]&r_1_addr[13]&r_0_addr[1],
r_2_addr[8]&r_1_addr[13]&r_0_addr[0],
r_2_addr[8]&r_1_addr[12]&r_0_addr[15],
r_2_addr[8]&r_1_addr[12]&r_0_addr[14],
r_2_addr[8]&r_1_addr[12]&r_0_addr[13],
r_2_addr[8]&r_1_addr[12]&r_0_addr[12],
r_2_addr[8]&r_1_addr[12]&r_0_addr[11],
r_2_addr[8]&r_1_addr[12]&r_0_addr[10],
r_2_addr[8]&r_1_addr[12]&r_0_addr[9],
r_2_addr[8]&r_1_addr[12]&r_0_addr[8],
r_2_addr[8]&r_1_addr[12]&r_0_addr[7],
r_2_addr[8]&r_1_addr[12]&r_0_addr[6],
r_2_addr[8]&r_1_addr[12]&r_0_addr[5],
r_2_addr[8]&r_1_addr[12]&r_0_addr[4],
r_2_addr[8]&r_1_addr[12]&r_0_addr[3],
r_2_addr[8]&r_1_addr[12]&r_0_addr[2],
r_2_addr[8]&r_1_addr[12]&r_0_addr[1],
r_2_addr[8]&r_1_addr[12]&r_0_addr[0],
r_2_addr[8]&r_1_addr[11]&r_0_addr[15],
r_2_addr[8]&r_1_addr[11]&r_0_addr[14],
r_2_addr[8]&r_1_addr[11]&r_0_addr[13],
r_2_addr[8]&r_1_addr[11]&r_0_addr[12],
r_2_addr[8]&r_1_addr[11]&r_0_addr[11],
r_2_addr[8]&r_1_addr[11]&r_0_addr[10],
r_2_addr[8]&r_1_addr[11]&r_0_addr[9],
r_2_addr[8]&r_1_addr[11]&r_0_addr[8],
r_2_addr[8]&r_1_addr[11]&r_0_addr[7],
r_2_addr[8]&r_1_addr[11]&r_0_addr[6],
r_2_addr[8]&r_1_addr[11]&r_0_addr[5],
r_2_addr[8]&r_1_addr[11]&r_0_addr[4],
r_2_addr[8]&r_1_addr[11]&r_0_addr[3],
r_2_addr[8]&r_1_addr[11]&r_0_addr[2],
r_2_addr[8]&r_1_addr[11]&r_0_addr[1],
r_2_addr[8]&r_1_addr[11]&r_0_addr[0],
r_2_addr[8]&r_1_addr[10]&r_0_addr[15],
r_2_addr[8]&r_1_addr[10]&r_0_addr[14],
r_2_addr[8]&r_1_addr[10]&r_0_addr[13],
r_2_addr[8]&r_1_addr[10]&r_0_addr[12],
r_2_addr[8]&r_1_addr[10]&r_0_addr[11],
r_2_addr[8]&r_1_addr[10]&r_0_addr[10],
r_2_addr[8]&r_1_addr[10]&r_0_addr[9],
r_2_addr[8]&r_1_addr[10]&r_0_addr[8],
r_2_addr[8]&r_1_addr[10]&r_0_addr[7],
r_2_addr[8]&r_1_addr[10]&r_0_addr[6],
r_2_addr[8]&r_1_addr[10]&r_0_addr[5],
r_2_addr[8]&r_1_addr[10]&r_0_addr[4],
r_2_addr[8]&r_1_addr[10]&r_0_addr[3],
r_2_addr[8]&r_1_addr[10]&r_0_addr[2],
r_2_addr[8]&r_1_addr[10]&r_0_addr[1],
r_2_addr[8]&r_1_addr[10]&r_0_addr[0],
r_2_addr[8]&r_1_addr[9]&r_0_addr[15],
r_2_addr[8]&r_1_addr[9]&r_0_addr[14],
r_2_addr[8]&r_1_addr[9]&r_0_addr[13],
r_2_addr[8]&r_1_addr[9]&r_0_addr[12],
r_2_addr[8]&r_1_addr[9]&r_0_addr[11],
r_2_addr[8]&r_1_addr[9]&r_0_addr[10],
r_2_addr[8]&r_1_addr[9]&r_0_addr[9],
r_2_addr[8]&r_1_addr[9]&r_0_addr[8],
r_2_addr[8]&r_1_addr[9]&r_0_addr[7],
r_2_addr[8]&r_1_addr[9]&r_0_addr[6],
r_2_addr[8]&r_1_addr[9]&r_0_addr[5],
r_2_addr[8]&r_1_addr[9]&r_0_addr[4],
r_2_addr[8]&r_1_addr[9]&r_0_addr[3],
r_2_addr[8]&r_1_addr[9]&r_0_addr[2],
r_2_addr[8]&r_1_addr[9]&r_0_addr[1],
r_2_addr[8]&r_1_addr[9]&r_0_addr[0],
r_2_addr[8]&r_1_addr[8]&r_0_addr[15],
r_2_addr[8]&r_1_addr[8]&r_0_addr[14],
r_2_addr[8]&r_1_addr[8]&r_0_addr[13],
r_2_addr[8]&r_1_addr[8]&r_0_addr[12],
r_2_addr[8]&r_1_addr[8]&r_0_addr[11],
r_2_addr[8]&r_1_addr[8]&r_0_addr[10],
r_2_addr[8]&r_1_addr[8]&r_0_addr[9],
r_2_addr[8]&r_1_addr[8]&r_0_addr[8],
r_2_addr[8]&r_1_addr[8]&r_0_addr[7],
r_2_addr[8]&r_1_addr[8]&r_0_addr[6],
r_2_addr[8]&r_1_addr[8]&r_0_addr[5],
r_2_addr[8]&r_1_addr[8]&r_0_addr[4],
r_2_addr[8]&r_1_addr[8]&r_0_addr[3],
r_2_addr[8]&r_1_addr[8]&r_0_addr[2],
r_2_addr[8]&r_1_addr[8]&r_0_addr[1],
r_2_addr[8]&r_1_addr[8]&r_0_addr[0],
r_2_addr[8]&r_1_addr[7]&r_0_addr[15],
r_2_addr[8]&r_1_addr[7]&r_0_addr[14],
r_2_addr[8]&r_1_addr[7]&r_0_addr[13],
r_2_addr[8]&r_1_addr[7]&r_0_addr[12],
r_2_addr[8]&r_1_addr[7]&r_0_addr[11],
r_2_addr[8]&r_1_addr[7]&r_0_addr[10],
r_2_addr[8]&r_1_addr[7]&r_0_addr[9],
r_2_addr[8]&r_1_addr[7]&r_0_addr[8],
r_2_addr[8]&r_1_addr[7]&r_0_addr[7],
r_2_addr[8]&r_1_addr[7]&r_0_addr[6],
r_2_addr[8]&r_1_addr[7]&r_0_addr[5],
r_2_addr[8]&r_1_addr[7]&r_0_addr[4],
r_2_addr[8]&r_1_addr[7]&r_0_addr[3],
r_2_addr[8]&r_1_addr[7]&r_0_addr[2],
r_2_addr[8]&r_1_addr[7]&r_0_addr[1],
r_2_addr[8]&r_1_addr[7]&r_0_addr[0],
r_2_addr[8]&r_1_addr[6]&r_0_addr[15],
r_2_addr[8]&r_1_addr[6]&r_0_addr[14],
r_2_addr[8]&r_1_addr[6]&r_0_addr[13],
r_2_addr[8]&r_1_addr[6]&r_0_addr[12],
r_2_addr[8]&r_1_addr[6]&r_0_addr[11],
r_2_addr[8]&r_1_addr[6]&r_0_addr[10],
r_2_addr[8]&r_1_addr[6]&r_0_addr[9],
r_2_addr[8]&r_1_addr[6]&r_0_addr[8],
r_2_addr[8]&r_1_addr[6]&r_0_addr[7],
r_2_addr[8]&r_1_addr[6]&r_0_addr[6],
r_2_addr[8]&r_1_addr[6]&r_0_addr[5],
r_2_addr[8]&r_1_addr[6]&r_0_addr[4],
r_2_addr[8]&r_1_addr[6]&r_0_addr[3],
r_2_addr[8]&r_1_addr[6]&r_0_addr[2],
r_2_addr[8]&r_1_addr[6]&r_0_addr[1],
r_2_addr[8]&r_1_addr[6]&r_0_addr[0],
r_2_addr[8]&r_1_addr[5]&r_0_addr[15],
r_2_addr[8]&r_1_addr[5]&r_0_addr[14],
r_2_addr[8]&r_1_addr[5]&r_0_addr[13],
r_2_addr[8]&r_1_addr[5]&r_0_addr[12],
r_2_addr[8]&r_1_addr[5]&r_0_addr[11],
r_2_addr[8]&r_1_addr[5]&r_0_addr[10],
r_2_addr[8]&r_1_addr[5]&r_0_addr[9],
r_2_addr[8]&r_1_addr[5]&r_0_addr[8],
r_2_addr[8]&r_1_addr[5]&r_0_addr[7],
r_2_addr[8]&r_1_addr[5]&r_0_addr[6],
r_2_addr[8]&r_1_addr[5]&r_0_addr[5],
r_2_addr[8]&r_1_addr[5]&r_0_addr[4],
r_2_addr[8]&r_1_addr[5]&r_0_addr[3],
r_2_addr[8]&r_1_addr[5]&r_0_addr[2],
r_2_addr[8]&r_1_addr[5]&r_0_addr[1],
r_2_addr[8]&r_1_addr[5]&r_0_addr[0],
r_2_addr[8]&r_1_addr[4]&r_0_addr[15],
r_2_addr[8]&r_1_addr[4]&r_0_addr[14],
r_2_addr[8]&r_1_addr[4]&r_0_addr[13],
r_2_addr[8]&r_1_addr[4]&r_0_addr[12],
r_2_addr[8]&r_1_addr[4]&r_0_addr[11],
r_2_addr[8]&r_1_addr[4]&r_0_addr[10],
r_2_addr[8]&r_1_addr[4]&r_0_addr[9],
r_2_addr[8]&r_1_addr[4]&r_0_addr[8],
r_2_addr[8]&r_1_addr[4]&r_0_addr[7],
r_2_addr[8]&r_1_addr[4]&r_0_addr[6],
r_2_addr[8]&r_1_addr[4]&r_0_addr[5],
r_2_addr[8]&r_1_addr[4]&r_0_addr[4],
r_2_addr[8]&r_1_addr[4]&r_0_addr[3],
r_2_addr[8]&r_1_addr[4]&r_0_addr[2],
r_2_addr[8]&r_1_addr[4]&r_0_addr[1],
r_2_addr[8]&r_1_addr[4]&r_0_addr[0],
r_2_addr[8]&r_1_addr[3]&r_0_addr[15],
r_2_addr[8]&r_1_addr[3]&r_0_addr[14],
r_2_addr[8]&r_1_addr[3]&r_0_addr[13],
r_2_addr[8]&r_1_addr[3]&r_0_addr[12],
r_2_addr[8]&r_1_addr[3]&r_0_addr[11],
r_2_addr[8]&r_1_addr[3]&r_0_addr[10],
r_2_addr[8]&r_1_addr[3]&r_0_addr[9],
r_2_addr[8]&r_1_addr[3]&r_0_addr[8],
r_2_addr[8]&r_1_addr[3]&r_0_addr[7],
r_2_addr[8]&r_1_addr[3]&r_0_addr[6],
r_2_addr[8]&r_1_addr[3]&r_0_addr[5],
r_2_addr[8]&r_1_addr[3]&r_0_addr[4],
r_2_addr[8]&r_1_addr[3]&r_0_addr[3],
r_2_addr[8]&r_1_addr[3]&r_0_addr[2],
r_2_addr[8]&r_1_addr[3]&r_0_addr[1],
r_2_addr[8]&r_1_addr[3]&r_0_addr[0],
r_2_addr[8]&r_1_addr[2]&r_0_addr[15],
r_2_addr[8]&r_1_addr[2]&r_0_addr[14],
r_2_addr[8]&r_1_addr[2]&r_0_addr[13],
r_2_addr[8]&r_1_addr[2]&r_0_addr[12],
r_2_addr[8]&r_1_addr[2]&r_0_addr[11],
r_2_addr[8]&r_1_addr[2]&r_0_addr[10],
r_2_addr[8]&r_1_addr[2]&r_0_addr[9],
r_2_addr[8]&r_1_addr[2]&r_0_addr[8],
r_2_addr[8]&r_1_addr[2]&r_0_addr[7],
r_2_addr[8]&r_1_addr[2]&r_0_addr[6],
r_2_addr[8]&r_1_addr[2]&r_0_addr[5],
r_2_addr[8]&r_1_addr[2]&r_0_addr[4],
r_2_addr[8]&r_1_addr[2]&r_0_addr[3],
r_2_addr[8]&r_1_addr[2]&r_0_addr[2],
r_2_addr[8]&r_1_addr[2]&r_0_addr[1],
r_2_addr[8]&r_1_addr[2]&r_0_addr[0],
r_2_addr[8]&r_1_addr[1]&r_0_addr[15],
r_2_addr[8]&r_1_addr[1]&r_0_addr[14],
r_2_addr[8]&r_1_addr[1]&r_0_addr[13],
r_2_addr[8]&r_1_addr[1]&r_0_addr[12],
r_2_addr[8]&r_1_addr[1]&r_0_addr[11],
r_2_addr[8]&r_1_addr[1]&r_0_addr[10],
r_2_addr[8]&r_1_addr[1]&r_0_addr[9],
r_2_addr[8]&r_1_addr[1]&r_0_addr[8],
r_2_addr[8]&r_1_addr[1]&r_0_addr[7],
r_2_addr[8]&r_1_addr[1]&r_0_addr[6],
r_2_addr[8]&r_1_addr[1]&r_0_addr[5],
r_2_addr[8]&r_1_addr[1]&r_0_addr[4],
r_2_addr[8]&r_1_addr[1]&r_0_addr[3],
r_2_addr[8]&r_1_addr[1]&r_0_addr[2],
r_2_addr[8]&r_1_addr[1]&r_0_addr[1],
r_2_addr[8]&r_1_addr[1]&r_0_addr[0],
r_2_addr[8]&r_1_addr[0]&r_0_addr[15],
r_2_addr[8]&r_1_addr[0]&r_0_addr[14],
r_2_addr[8]&r_1_addr[0]&r_0_addr[13],
r_2_addr[8]&r_1_addr[0]&r_0_addr[12],
r_2_addr[8]&r_1_addr[0]&r_0_addr[11],
r_2_addr[8]&r_1_addr[0]&r_0_addr[10],
r_2_addr[8]&r_1_addr[0]&r_0_addr[9],
r_2_addr[8]&r_1_addr[0]&r_0_addr[8],
r_2_addr[8]&r_1_addr[0]&r_0_addr[7],
r_2_addr[8]&r_1_addr[0]&r_0_addr[6],
r_2_addr[8]&r_1_addr[0]&r_0_addr[5],
r_2_addr[8]&r_1_addr[0]&r_0_addr[4],
r_2_addr[8]&r_1_addr[0]&r_0_addr[3],
r_2_addr[8]&r_1_addr[0]&r_0_addr[2],
r_2_addr[8]&r_1_addr[0]&r_0_addr[1],
r_2_addr[8]&r_1_addr[0]&r_0_addr[0],
r_2_addr[7]&r_1_addr[15]&r_0_addr[15],
r_2_addr[7]&r_1_addr[15]&r_0_addr[14],
r_2_addr[7]&r_1_addr[15]&r_0_addr[13],
r_2_addr[7]&r_1_addr[15]&r_0_addr[12],
r_2_addr[7]&r_1_addr[15]&r_0_addr[11],
r_2_addr[7]&r_1_addr[15]&r_0_addr[10],
r_2_addr[7]&r_1_addr[15]&r_0_addr[9],
r_2_addr[7]&r_1_addr[15]&r_0_addr[8],
r_2_addr[7]&r_1_addr[15]&r_0_addr[7],
r_2_addr[7]&r_1_addr[15]&r_0_addr[6],
r_2_addr[7]&r_1_addr[15]&r_0_addr[5],
r_2_addr[7]&r_1_addr[15]&r_0_addr[4],
r_2_addr[7]&r_1_addr[15]&r_0_addr[3],
r_2_addr[7]&r_1_addr[15]&r_0_addr[2],
r_2_addr[7]&r_1_addr[15]&r_0_addr[1],
r_2_addr[7]&r_1_addr[15]&r_0_addr[0],
r_2_addr[7]&r_1_addr[14]&r_0_addr[15],
r_2_addr[7]&r_1_addr[14]&r_0_addr[14],
r_2_addr[7]&r_1_addr[14]&r_0_addr[13],
r_2_addr[7]&r_1_addr[14]&r_0_addr[12],
r_2_addr[7]&r_1_addr[14]&r_0_addr[11],
r_2_addr[7]&r_1_addr[14]&r_0_addr[10],
r_2_addr[7]&r_1_addr[14]&r_0_addr[9],
r_2_addr[7]&r_1_addr[14]&r_0_addr[8],
r_2_addr[7]&r_1_addr[14]&r_0_addr[7],
r_2_addr[7]&r_1_addr[14]&r_0_addr[6],
r_2_addr[7]&r_1_addr[14]&r_0_addr[5],
r_2_addr[7]&r_1_addr[14]&r_0_addr[4],
r_2_addr[7]&r_1_addr[14]&r_0_addr[3],
r_2_addr[7]&r_1_addr[14]&r_0_addr[2],
r_2_addr[7]&r_1_addr[14]&r_0_addr[1],
r_2_addr[7]&r_1_addr[14]&r_0_addr[0],
r_2_addr[7]&r_1_addr[13]&r_0_addr[15],
r_2_addr[7]&r_1_addr[13]&r_0_addr[14],
r_2_addr[7]&r_1_addr[13]&r_0_addr[13],
r_2_addr[7]&r_1_addr[13]&r_0_addr[12],
r_2_addr[7]&r_1_addr[13]&r_0_addr[11],
r_2_addr[7]&r_1_addr[13]&r_0_addr[10],
r_2_addr[7]&r_1_addr[13]&r_0_addr[9],
r_2_addr[7]&r_1_addr[13]&r_0_addr[8],
r_2_addr[7]&r_1_addr[13]&r_0_addr[7],
r_2_addr[7]&r_1_addr[13]&r_0_addr[6],
r_2_addr[7]&r_1_addr[13]&r_0_addr[5],
r_2_addr[7]&r_1_addr[13]&r_0_addr[4],
r_2_addr[7]&r_1_addr[13]&r_0_addr[3],
r_2_addr[7]&r_1_addr[13]&r_0_addr[2],
r_2_addr[7]&r_1_addr[13]&r_0_addr[1],
r_2_addr[7]&r_1_addr[13]&r_0_addr[0],
r_2_addr[7]&r_1_addr[12]&r_0_addr[15],
r_2_addr[7]&r_1_addr[12]&r_0_addr[14],
r_2_addr[7]&r_1_addr[12]&r_0_addr[13],
r_2_addr[7]&r_1_addr[12]&r_0_addr[12],
r_2_addr[7]&r_1_addr[12]&r_0_addr[11],
r_2_addr[7]&r_1_addr[12]&r_0_addr[10],
r_2_addr[7]&r_1_addr[12]&r_0_addr[9],
r_2_addr[7]&r_1_addr[12]&r_0_addr[8],
r_2_addr[7]&r_1_addr[12]&r_0_addr[7],
r_2_addr[7]&r_1_addr[12]&r_0_addr[6],
r_2_addr[7]&r_1_addr[12]&r_0_addr[5],
r_2_addr[7]&r_1_addr[12]&r_0_addr[4],
r_2_addr[7]&r_1_addr[12]&r_0_addr[3],
r_2_addr[7]&r_1_addr[12]&r_0_addr[2],
r_2_addr[7]&r_1_addr[12]&r_0_addr[1],
r_2_addr[7]&r_1_addr[12]&r_0_addr[0],
r_2_addr[7]&r_1_addr[11]&r_0_addr[15],
r_2_addr[7]&r_1_addr[11]&r_0_addr[14],
r_2_addr[7]&r_1_addr[11]&r_0_addr[13],
r_2_addr[7]&r_1_addr[11]&r_0_addr[12],
r_2_addr[7]&r_1_addr[11]&r_0_addr[11],
r_2_addr[7]&r_1_addr[11]&r_0_addr[10],
r_2_addr[7]&r_1_addr[11]&r_0_addr[9],
r_2_addr[7]&r_1_addr[11]&r_0_addr[8],
r_2_addr[7]&r_1_addr[11]&r_0_addr[7],
r_2_addr[7]&r_1_addr[11]&r_0_addr[6],
r_2_addr[7]&r_1_addr[11]&r_0_addr[5],
r_2_addr[7]&r_1_addr[11]&r_0_addr[4],
r_2_addr[7]&r_1_addr[11]&r_0_addr[3],
r_2_addr[7]&r_1_addr[11]&r_0_addr[2],
r_2_addr[7]&r_1_addr[11]&r_0_addr[1],
r_2_addr[7]&r_1_addr[11]&r_0_addr[0],
r_2_addr[7]&r_1_addr[10]&r_0_addr[15],
r_2_addr[7]&r_1_addr[10]&r_0_addr[14],
r_2_addr[7]&r_1_addr[10]&r_0_addr[13],
r_2_addr[7]&r_1_addr[10]&r_0_addr[12],
r_2_addr[7]&r_1_addr[10]&r_0_addr[11],
r_2_addr[7]&r_1_addr[10]&r_0_addr[10],
r_2_addr[7]&r_1_addr[10]&r_0_addr[9],
r_2_addr[7]&r_1_addr[10]&r_0_addr[8],
r_2_addr[7]&r_1_addr[10]&r_0_addr[7],
r_2_addr[7]&r_1_addr[10]&r_0_addr[6],
r_2_addr[7]&r_1_addr[10]&r_0_addr[5],
r_2_addr[7]&r_1_addr[10]&r_0_addr[4],
r_2_addr[7]&r_1_addr[10]&r_0_addr[3],
r_2_addr[7]&r_1_addr[10]&r_0_addr[2],
r_2_addr[7]&r_1_addr[10]&r_0_addr[1],
r_2_addr[7]&r_1_addr[10]&r_0_addr[0],
r_2_addr[7]&r_1_addr[9]&r_0_addr[15],
r_2_addr[7]&r_1_addr[9]&r_0_addr[14],
r_2_addr[7]&r_1_addr[9]&r_0_addr[13],
r_2_addr[7]&r_1_addr[9]&r_0_addr[12],
r_2_addr[7]&r_1_addr[9]&r_0_addr[11],
r_2_addr[7]&r_1_addr[9]&r_0_addr[10],
r_2_addr[7]&r_1_addr[9]&r_0_addr[9],
r_2_addr[7]&r_1_addr[9]&r_0_addr[8],
r_2_addr[7]&r_1_addr[9]&r_0_addr[7],
r_2_addr[7]&r_1_addr[9]&r_0_addr[6],
r_2_addr[7]&r_1_addr[9]&r_0_addr[5],
r_2_addr[7]&r_1_addr[9]&r_0_addr[4],
r_2_addr[7]&r_1_addr[9]&r_0_addr[3],
r_2_addr[7]&r_1_addr[9]&r_0_addr[2],
r_2_addr[7]&r_1_addr[9]&r_0_addr[1],
r_2_addr[7]&r_1_addr[9]&r_0_addr[0],
r_2_addr[7]&r_1_addr[8]&r_0_addr[15],
r_2_addr[7]&r_1_addr[8]&r_0_addr[14],
r_2_addr[7]&r_1_addr[8]&r_0_addr[13],
r_2_addr[7]&r_1_addr[8]&r_0_addr[12],
r_2_addr[7]&r_1_addr[8]&r_0_addr[11],
r_2_addr[7]&r_1_addr[8]&r_0_addr[10],
r_2_addr[7]&r_1_addr[8]&r_0_addr[9],
r_2_addr[7]&r_1_addr[8]&r_0_addr[8],
r_2_addr[7]&r_1_addr[8]&r_0_addr[7],
r_2_addr[7]&r_1_addr[8]&r_0_addr[6],
r_2_addr[7]&r_1_addr[8]&r_0_addr[5],
r_2_addr[7]&r_1_addr[8]&r_0_addr[4],
r_2_addr[7]&r_1_addr[8]&r_0_addr[3],
r_2_addr[7]&r_1_addr[8]&r_0_addr[2],
r_2_addr[7]&r_1_addr[8]&r_0_addr[1],
r_2_addr[7]&r_1_addr[8]&r_0_addr[0],
r_2_addr[7]&r_1_addr[7]&r_0_addr[15],
r_2_addr[7]&r_1_addr[7]&r_0_addr[14],
r_2_addr[7]&r_1_addr[7]&r_0_addr[13],
r_2_addr[7]&r_1_addr[7]&r_0_addr[12],
r_2_addr[7]&r_1_addr[7]&r_0_addr[11],
r_2_addr[7]&r_1_addr[7]&r_0_addr[10],
r_2_addr[7]&r_1_addr[7]&r_0_addr[9],
r_2_addr[7]&r_1_addr[7]&r_0_addr[8],
r_2_addr[7]&r_1_addr[7]&r_0_addr[7],
r_2_addr[7]&r_1_addr[7]&r_0_addr[6],
r_2_addr[7]&r_1_addr[7]&r_0_addr[5],
r_2_addr[7]&r_1_addr[7]&r_0_addr[4],
r_2_addr[7]&r_1_addr[7]&r_0_addr[3],
r_2_addr[7]&r_1_addr[7]&r_0_addr[2],
r_2_addr[7]&r_1_addr[7]&r_0_addr[1],
r_2_addr[7]&r_1_addr[7]&r_0_addr[0],
r_2_addr[7]&r_1_addr[6]&r_0_addr[15],
r_2_addr[7]&r_1_addr[6]&r_0_addr[14],
r_2_addr[7]&r_1_addr[6]&r_0_addr[13],
r_2_addr[7]&r_1_addr[6]&r_0_addr[12],
r_2_addr[7]&r_1_addr[6]&r_0_addr[11],
r_2_addr[7]&r_1_addr[6]&r_0_addr[10],
r_2_addr[7]&r_1_addr[6]&r_0_addr[9],
r_2_addr[7]&r_1_addr[6]&r_0_addr[8],
r_2_addr[7]&r_1_addr[6]&r_0_addr[7],
r_2_addr[7]&r_1_addr[6]&r_0_addr[6],
r_2_addr[7]&r_1_addr[6]&r_0_addr[5],
r_2_addr[7]&r_1_addr[6]&r_0_addr[4],
r_2_addr[7]&r_1_addr[6]&r_0_addr[3],
r_2_addr[7]&r_1_addr[6]&r_0_addr[2],
r_2_addr[7]&r_1_addr[6]&r_0_addr[1],
r_2_addr[7]&r_1_addr[6]&r_0_addr[0],
r_2_addr[7]&r_1_addr[5]&r_0_addr[15],
r_2_addr[7]&r_1_addr[5]&r_0_addr[14],
r_2_addr[7]&r_1_addr[5]&r_0_addr[13],
r_2_addr[7]&r_1_addr[5]&r_0_addr[12],
r_2_addr[7]&r_1_addr[5]&r_0_addr[11],
r_2_addr[7]&r_1_addr[5]&r_0_addr[10],
r_2_addr[7]&r_1_addr[5]&r_0_addr[9],
r_2_addr[7]&r_1_addr[5]&r_0_addr[8],
r_2_addr[7]&r_1_addr[5]&r_0_addr[7],
r_2_addr[7]&r_1_addr[5]&r_0_addr[6],
r_2_addr[7]&r_1_addr[5]&r_0_addr[5],
r_2_addr[7]&r_1_addr[5]&r_0_addr[4],
r_2_addr[7]&r_1_addr[5]&r_0_addr[3],
r_2_addr[7]&r_1_addr[5]&r_0_addr[2],
r_2_addr[7]&r_1_addr[5]&r_0_addr[1],
r_2_addr[7]&r_1_addr[5]&r_0_addr[0],
r_2_addr[7]&r_1_addr[4]&r_0_addr[15],
r_2_addr[7]&r_1_addr[4]&r_0_addr[14],
r_2_addr[7]&r_1_addr[4]&r_0_addr[13],
r_2_addr[7]&r_1_addr[4]&r_0_addr[12],
r_2_addr[7]&r_1_addr[4]&r_0_addr[11],
r_2_addr[7]&r_1_addr[4]&r_0_addr[10],
r_2_addr[7]&r_1_addr[4]&r_0_addr[9],
r_2_addr[7]&r_1_addr[4]&r_0_addr[8],
r_2_addr[7]&r_1_addr[4]&r_0_addr[7],
r_2_addr[7]&r_1_addr[4]&r_0_addr[6],
r_2_addr[7]&r_1_addr[4]&r_0_addr[5],
r_2_addr[7]&r_1_addr[4]&r_0_addr[4],
r_2_addr[7]&r_1_addr[4]&r_0_addr[3],
r_2_addr[7]&r_1_addr[4]&r_0_addr[2],
r_2_addr[7]&r_1_addr[4]&r_0_addr[1],
r_2_addr[7]&r_1_addr[4]&r_0_addr[0],
r_2_addr[7]&r_1_addr[3]&r_0_addr[15],
r_2_addr[7]&r_1_addr[3]&r_0_addr[14],
r_2_addr[7]&r_1_addr[3]&r_0_addr[13],
r_2_addr[7]&r_1_addr[3]&r_0_addr[12],
r_2_addr[7]&r_1_addr[3]&r_0_addr[11],
r_2_addr[7]&r_1_addr[3]&r_0_addr[10],
r_2_addr[7]&r_1_addr[3]&r_0_addr[9],
r_2_addr[7]&r_1_addr[3]&r_0_addr[8],
r_2_addr[7]&r_1_addr[3]&r_0_addr[7],
r_2_addr[7]&r_1_addr[3]&r_0_addr[6],
r_2_addr[7]&r_1_addr[3]&r_0_addr[5],
r_2_addr[7]&r_1_addr[3]&r_0_addr[4],
r_2_addr[7]&r_1_addr[3]&r_0_addr[3],
r_2_addr[7]&r_1_addr[3]&r_0_addr[2],
r_2_addr[7]&r_1_addr[3]&r_0_addr[1],
r_2_addr[7]&r_1_addr[3]&r_0_addr[0],
r_2_addr[7]&r_1_addr[2]&r_0_addr[15],
r_2_addr[7]&r_1_addr[2]&r_0_addr[14],
r_2_addr[7]&r_1_addr[2]&r_0_addr[13],
r_2_addr[7]&r_1_addr[2]&r_0_addr[12],
r_2_addr[7]&r_1_addr[2]&r_0_addr[11],
r_2_addr[7]&r_1_addr[2]&r_0_addr[10],
r_2_addr[7]&r_1_addr[2]&r_0_addr[9],
r_2_addr[7]&r_1_addr[2]&r_0_addr[8],
r_2_addr[7]&r_1_addr[2]&r_0_addr[7],
r_2_addr[7]&r_1_addr[2]&r_0_addr[6],
r_2_addr[7]&r_1_addr[2]&r_0_addr[5],
r_2_addr[7]&r_1_addr[2]&r_0_addr[4],
r_2_addr[7]&r_1_addr[2]&r_0_addr[3],
r_2_addr[7]&r_1_addr[2]&r_0_addr[2],
r_2_addr[7]&r_1_addr[2]&r_0_addr[1],
r_2_addr[7]&r_1_addr[2]&r_0_addr[0],
r_2_addr[7]&r_1_addr[1]&r_0_addr[15],
r_2_addr[7]&r_1_addr[1]&r_0_addr[14],
r_2_addr[7]&r_1_addr[1]&r_0_addr[13],
r_2_addr[7]&r_1_addr[1]&r_0_addr[12],
r_2_addr[7]&r_1_addr[1]&r_0_addr[11],
r_2_addr[7]&r_1_addr[1]&r_0_addr[10],
r_2_addr[7]&r_1_addr[1]&r_0_addr[9],
r_2_addr[7]&r_1_addr[1]&r_0_addr[8],
r_2_addr[7]&r_1_addr[1]&r_0_addr[7],
r_2_addr[7]&r_1_addr[1]&r_0_addr[6],
r_2_addr[7]&r_1_addr[1]&r_0_addr[5],
r_2_addr[7]&r_1_addr[1]&r_0_addr[4],
r_2_addr[7]&r_1_addr[1]&r_0_addr[3],
r_2_addr[7]&r_1_addr[1]&r_0_addr[2],
r_2_addr[7]&r_1_addr[1]&r_0_addr[1],
r_2_addr[7]&r_1_addr[1]&r_0_addr[0],
r_2_addr[7]&r_1_addr[0]&r_0_addr[15],
r_2_addr[7]&r_1_addr[0]&r_0_addr[14],
r_2_addr[7]&r_1_addr[0]&r_0_addr[13],
r_2_addr[7]&r_1_addr[0]&r_0_addr[12],
r_2_addr[7]&r_1_addr[0]&r_0_addr[11],
r_2_addr[7]&r_1_addr[0]&r_0_addr[10],
r_2_addr[7]&r_1_addr[0]&r_0_addr[9],
r_2_addr[7]&r_1_addr[0]&r_0_addr[8],
r_2_addr[7]&r_1_addr[0]&r_0_addr[7],
r_2_addr[7]&r_1_addr[0]&r_0_addr[6],
r_2_addr[7]&r_1_addr[0]&r_0_addr[5],
r_2_addr[7]&r_1_addr[0]&r_0_addr[4],
r_2_addr[7]&r_1_addr[0]&r_0_addr[3],
r_2_addr[7]&r_1_addr[0]&r_0_addr[2],
r_2_addr[7]&r_1_addr[0]&r_0_addr[1],
r_2_addr[7]&r_1_addr[0]&r_0_addr[0],
r_2_addr[6]&r_1_addr[15]&r_0_addr[15],
r_2_addr[6]&r_1_addr[15]&r_0_addr[14],
r_2_addr[6]&r_1_addr[15]&r_0_addr[13],
r_2_addr[6]&r_1_addr[15]&r_0_addr[12],
r_2_addr[6]&r_1_addr[15]&r_0_addr[11],
r_2_addr[6]&r_1_addr[15]&r_0_addr[10],
r_2_addr[6]&r_1_addr[15]&r_0_addr[9],
r_2_addr[6]&r_1_addr[15]&r_0_addr[8],
r_2_addr[6]&r_1_addr[15]&r_0_addr[7],
r_2_addr[6]&r_1_addr[15]&r_0_addr[6],
r_2_addr[6]&r_1_addr[15]&r_0_addr[5],
r_2_addr[6]&r_1_addr[15]&r_0_addr[4],
r_2_addr[6]&r_1_addr[15]&r_0_addr[3],
r_2_addr[6]&r_1_addr[15]&r_0_addr[2],
r_2_addr[6]&r_1_addr[15]&r_0_addr[1],
r_2_addr[6]&r_1_addr[15]&r_0_addr[0],
r_2_addr[6]&r_1_addr[14]&r_0_addr[15],
r_2_addr[6]&r_1_addr[14]&r_0_addr[14],
r_2_addr[6]&r_1_addr[14]&r_0_addr[13],
r_2_addr[6]&r_1_addr[14]&r_0_addr[12],
r_2_addr[6]&r_1_addr[14]&r_0_addr[11],
r_2_addr[6]&r_1_addr[14]&r_0_addr[10],
r_2_addr[6]&r_1_addr[14]&r_0_addr[9],
r_2_addr[6]&r_1_addr[14]&r_0_addr[8],
r_2_addr[6]&r_1_addr[14]&r_0_addr[7],
r_2_addr[6]&r_1_addr[14]&r_0_addr[6],
r_2_addr[6]&r_1_addr[14]&r_0_addr[5],
r_2_addr[6]&r_1_addr[14]&r_0_addr[4],
r_2_addr[6]&r_1_addr[14]&r_0_addr[3],
r_2_addr[6]&r_1_addr[14]&r_0_addr[2],
r_2_addr[6]&r_1_addr[14]&r_0_addr[1],
r_2_addr[6]&r_1_addr[14]&r_0_addr[0],
r_2_addr[6]&r_1_addr[13]&r_0_addr[15],
r_2_addr[6]&r_1_addr[13]&r_0_addr[14],
r_2_addr[6]&r_1_addr[13]&r_0_addr[13],
r_2_addr[6]&r_1_addr[13]&r_0_addr[12],
r_2_addr[6]&r_1_addr[13]&r_0_addr[11],
r_2_addr[6]&r_1_addr[13]&r_0_addr[10],
r_2_addr[6]&r_1_addr[13]&r_0_addr[9],
r_2_addr[6]&r_1_addr[13]&r_0_addr[8],
r_2_addr[6]&r_1_addr[13]&r_0_addr[7],
r_2_addr[6]&r_1_addr[13]&r_0_addr[6],
r_2_addr[6]&r_1_addr[13]&r_0_addr[5],
r_2_addr[6]&r_1_addr[13]&r_0_addr[4],
r_2_addr[6]&r_1_addr[13]&r_0_addr[3],
r_2_addr[6]&r_1_addr[13]&r_0_addr[2],
r_2_addr[6]&r_1_addr[13]&r_0_addr[1],
r_2_addr[6]&r_1_addr[13]&r_0_addr[0],
r_2_addr[6]&r_1_addr[12]&r_0_addr[15],
r_2_addr[6]&r_1_addr[12]&r_0_addr[14],
r_2_addr[6]&r_1_addr[12]&r_0_addr[13],
r_2_addr[6]&r_1_addr[12]&r_0_addr[12],
r_2_addr[6]&r_1_addr[12]&r_0_addr[11],
r_2_addr[6]&r_1_addr[12]&r_0_addr[10],
r_2_addr[6]&r_1_addr[12]&r_0_addr[9],
r_2_addr[6]&r_1_addr[12]&r_0_addr[8],
r_2_addr[6]&r_1_addr[12]&r_0_addr[7],
r_2_addr[6]&r_1_addr[12]&r_0_addr[6],
r_2_addr[6]&r_1_addr[12]&r_0_addr[5],
r_2_addr[6]&r_1_addr[12]&r_0_addr[4],
r_2_addr[6]&r_1_addr[12]&r_0_addr[3],
r_2_addr[6]&r_1_addr[12]&r_0_addr[2],
r_2_addr[6]&r_1_addr[12]&r_0_addr[1],
r_2_addr[6]&r_1_addr[12]&r_0_addr[0],
r_2_addr[6]&r_1_addr[11]&r_0_addr[15],
r_2_addr[6]&r_1_addr[11]&r_0_addr[14],
r_2_addr[6]&r_1_addr[11]&r_0_addr[13],
r_2_addr[6]&r_1_addr[11]&r_0_addr[12],
r_2_addr[6]&r_1_addr[11]&r_0_addr[11],
r_2_addr[6]&r_1_addr[11]&r_0_addr[10],
r_2_addr[6]&r_1_addr[11]&r_0_addr[9],
r_2_addr[6]&r_1_addr[11]&r_0_addr[8],
r_2_addr[6]&r_1_addr[11]&r_0_addr[7],
r_2_addr[6]&r_1_addr[11]&r_0_addr[6],
r_2_addr[6]&r_1_addr[11]&r_0_addr[5],
r_2_addr[6]&r_1_addr[11]&r_0_addr[4],
r_2_addr[6]&r_1_addr[11]&r_0_addr[3],
r_2_addr[6]&r_1_addr[11]&r_0_addr[2],
r_2_addr[6]&r_1_addr[11]&r_0_addr[1],
r_2_addr[6]&r_1_addr[11]&r_0_addr[0],
r_2_addr[6]&r_1_addr[10]&r_0_addr[15],
r_2_addr[6]&r_1_addr[10]&r_0_addr[14],
r_2_addr[6]&r_1_addr[10]&r_0_addr[13],
r_2_addr[6]&r_1_addr[10]&r_0_addr[12],
r_2_addr[6]&r_1_addr[10]&r_0_addr[11],
r_2_addr[6]&r_1_addr[10]&r_0_addr[10],
r_2_addr[6]&r_1_addr[10]&r_0_addr[9],
r_2_addr[6]&r_1_addr[10]&r_0_addr[8],
r_2_addr[6]&r_1_addr[10]&r_0_addr[7],
r_2_addr[6]&r_1_addr[10]&r_0_addr[6],
r_2_addr[6]&r_1_addr[10]&r_0_addr[5],
r_2_addr[6]&r_1_addr[10]&r_0_addr[4],
r_2_addr[6]&r_1_addr[10]&r_0_addr[3],
r_2_addr[6]&r_1_addr[10]&r_0_addr[2],
r_2_addr[6]&r_1_addr[10]&r_0_addr[1],
r_2_addr[6]&r_1_addr[10]&r_0_addr[0],
r_2_addr[6]&r_1_addr[9]&r_0_addr[15],
r_2_addr[6]&r_1_addr[9]&r_0_addr[14],
r_2_addr[6]&r_1_addr[9]&r_0_addr[13],
r_2_addr[6]&r_1_addr[9]&r_0_addr[12],
r_2_addr[6]&r_1_addr[9]&r_0_addr[11],
r_2_addr[6]&r_1_addr[9]&r_0_addr[10],
r_2_addr[6]&r_1_addr[9]&r_0_addr[9],
r_2_addr[6]&r_1_addr[9]&r_0_addr[8],
r_2_addr[6]&r_1_addr[9]&r_0_addr[7],
r_2_addr[6]&r_1_addr[9]&r_0_addr[6],
r_2_addr[6]&r_1_addr[9]&r_0_addr[5],
r_2_addr[6]&r_1_addr[9]&r_0_addr[4],
r_2_addr[6]&r_1_addr[9]&r_0_addr[3],
r_2_addr[6]&r_1_addr[9]&r_0_addr[2],
r_2_addr[6]&r_1_addr[9]&r_0_addr[1],
r_2_addr[6]&r_1_addr[9]&r_0_addr[0],
r_2_addr[6]&r_1_addr[8]&r_0_addr[15],
r_2_addr[6]&r_1_addr[8]&r_0_addr[14],
r_2_addr[6]&r_1_addr[8]&r_0_addr[13],
r_2_addr[6]&r_1_addr[8]&r_0_addr[12],
r_2_addr[6]&r_1_addr[8]&r_0_addr[11],
r_2_addr[6]&r_1_addr[8]&r_0_addr[10],
r_2_addr[6]&r_1_addr[8]&r_0_addr[9],
r_2_addr[6]&r_1_addr[8]&r_0_addr[8],
r_2_addr[6]&r_1_addr[8]&r_0_addr[7],
r_2_addr[6]&r_1_addr[8]&r_0_addr[6],
r_2_addr[6]&r_1_addr[8]&r_0_addr[5],
r_2_addr[6]&r_1_addr[8]&r_0_addr[4],
r_2_addr[6]&r_1_addr[8]&r_0_addr[3],
r_2_addr[6]&r_1_addr[8]&r_0_addr[2],
r_2_addr[6]&r_1_addr[8]&r_0_addr[1],
r_2_addr[6]&r_1_addr[8]&r_0_addr[0],
r_2_addr[6]&r_1_addr[7]&r_0_addr[15],
r_2_addr[6]&r_1_addr[7]&r_0_addr[14],
r_2_addr[6]&r_1_addr[7]&r_0_addr[13],
r_2_addr[6]&r_1_addr[7]&r_0_addr[12],
r_2_addr[6]&r_1_addr[7]&r_0_addr[11],
r_2_addr[6]&r_1_addr[7]&r_0_addr[10],
r_2_addr[6]&r_1_addr[7]&r_0_addr[9],
r_2_addr[6]&r_1_addr[7]&r_0_addr[8],
r_2_addr[6]&r_1_addr[7]&r_0_addr[7],
r_2_addr[6]&r_1_addr[7]&r_0_addr[6],
r_2_addr[6]&r_1_addr[7]&r_0_addr[5],
r_2_addr[6]&r_1_addr[7]&r_0_addr[4],
r_2_addr[6]&r_1_addr[7]&r_0_addr[3],
r_2_addr[6]&r_1_addr[7]&r_0_addr[2],
r_2_addr[6]&r_1_addr[7]&r_0_addr[1],
r_2_addr[6]&r_1_addr[7]&r_0_addr[0],
r_2_addr[6]&r_1_addr[6]&r_0_addr[15],
r_2_addr[6]&r_1_addr[6]&r_0_addr[14],
r_2_addr[6]&r_1_addr[6]&r_0_addr[13],
r_2_addr[6]&r_1_addr[6]&r_0_addr[12],
r_2_addr[6]&r_1_addr[6]&r_0_addr[11],
r_2_addr[6]&r_1_addr[6]&r_0_addr[10],
r_2_addr[6]&r_1_addr[6]&r_0_addr[9],
r_2_addr[6]&r_1_addr[6]&r_0_addr[8],
r_2_addr[6]&r_1_addr[6]&r_0_addr[7],
r_2_addr[6]&r_1_addr[6]&r_0_addr[6],
r_2_addr[6]&r_1_addr[6]&r_0_addr[5],
r_2_addr[6]&r_1_addr[6]&r_0_addr[4],
r_2_addr[6]&r_1_addr[6]&r_0_addr[3],
r_2_addr[6]&r_1_addr[6]&r_0_addr[2],
r_2_addr[6]&r_1_addr[6]&r_0_addr[1],
r_2_addr[6]&r_1_addr[6]&r_0_addr[0],
r_2_addr[6]&r_1_addr[5]&r_0_addr[15],
r_2_addr[6]&r_1_addr[5]&r_0_addr[14],
r_2_addr[6]&r_1_addr[5]&r_0_addr[13],
r_2_addr[6]&r_1_addr[5]&r_0_addr[12],
r_2_addr[6]&r_1_addr[5]&r_0_addr[11],
r_2_addr[6]&r_1_addr[5]&r_0_addr[10],
r_2_addr[6]&r_1_addr[5]&r_0_addr[9],
r_2_addr[6]&r_1_addr[5]&r_0_addr[8],
r_2_addr[6]&r_1_addr[5]&r_0_addr[7],
r_2_addr[6]&r_1_addr[5]&r_0_addr[6],
r_2_addr[6]&r_1_addr[5]&r_0_addr[5],
r_2_addr[6]&r_1_addr[5]&r_0_addr[4],
r_2_addr[6]&r_1_addr[5]&r_0_addr[3],
r_2_addr[6]&r_1_addr[5]&r_0_addr[2],
r_2_addr[6]&r_1_addr[5]&r_0_addr[1],
r_2_addr[6]&r_1_addr[5]&r_0_addr[0],
r_2_addr[6]&r_1_addr[4]&r_0_addr[15],
r_2_addr[6]&r_1_addr[4]&r_0_addr[14],
r_2_addr[6]&r_1_addr[4]&r_0_addr[13],
r_2_addr[6]&r_1_addr[4]&r_0_addr[12],
r_2_addr[6]&r_1_addr[4]&r_0_addr[11],
r_2_addr[6]&r_1_addr[4]&r_0_addr[10],
r_2_addr[6]&r_1_addr[4]&r_0_addr[9],
r_2_addr[6]&r_1_addr[4]&r_0_addr[8],
r_2_addr[6]&r_1_addr[4]&r_0_addr[7],
r_2_addr[6]&r_1_addr[4]&r_0_addr[6],
r_2_addr[6]&r_1_addr[4]&r_0_addr[5],
r_2_addr[6]&r_1_addr[4]&r_0_addr[4],
r_2_addr[6]&r_1_addr[4]&r_0_addr[3],
r_2_addr[6]&r_1_addr[4]&r_0_addr[2],
r_2_addr[6]&r_1_addr[4]&r_0_addr[1],
r_2_addr[6]&r_1_addr[4]&r_0_addr[0],
r_2_addr[6]&r_1_addr[3]&r_0_addr[15],
r_2_addr[6]&r_1_addr[3]&r_0_addr[14],
r_2_addr[6]&r_1_addr[3]&r_0_addr[13],
r_2_addr[6]&r_1_addr[3]&r_0_addr[12],
r_2_addr[6]&r_1_addr[3]&r_0_addr[11],
r_2_addr[6]&r_1_addr[3]&r_0_addr[10],
r_2_addr[6]&r_1_addr[3]&r_0_addr[9],
r_2_addr[6]&r_1_addr[3]&r_0_addr[8],
r_2_addr[6]&r_1_addr[3]&r_0_addr[7],
r_2_addr[6]&r_1_addr[3]&r_0_addr[6],
r_2_addr[6]&r_1_addr[3]&r_0_addr[5],
r_2_addr[6]&r_1_addr[3]&r_0_addr[4],
r_2_addr[6]&r_1_addr[3]&r_0_addr[3],
r_2_addr[6]&r_1_addr[3]&r_0_addr[2],
r_2_addr[6]&r_1_addr[3]&r_0_addr[1],
r_2_addr[6]&r_1_addr[3]&r_0_addr[0],
r_2_addr[6]&r_1_addr[2]&r_0_addr[15],
r_2_addr[6]&r_1_addr[2]&r_0_addr[14],
r_2_addr[6]&r_1_addr[2]&r_0_addr[13],
r_2_addr[6]&r_1_addr[2]&r_0_addr[12],
r_2_addr[6]&r_1_addr[2]&r_0_addr[11],
r_2_addr[6]&r_1_addr[2]&r_0_addr[10],
r_2_addr[6]&r_1_addr[2]&r_0_addr[9],
r_2_addr[6]&r_1_addr[2]&r_0_addr[8],
r_2_addr[6]&r_1_addr[2]&r_0_addr[7],
r_2_addr[6]&r_1_addr[2]&r_0_addr[6],
r_2_addr[6]&r_1_addr[2]&r_0_addr[5],
r_2_addr[6]&r_1_addr[2]&r_0_addr[4],
r_2_addr[6]&r_1_addr[2]&r_0_addr[3],
r_2_addr[6]&r_1_addr[2]&r_0_addr[2],
r_2_addr[6]&r_1_addr[2]&r_0_addr[1],
r_2_addr[6]&r_1_addr[2]&r_0_addr[0],
r_2_addr[6]&r_1_addr[1]&r_0_addr[15],
r_2_addr[6]&r_1_addr[1]&r_0_addr[14],
r_2_addr[6]&r_1_addr[1]&r_0_addr[13],
r_2_addr[6]&r_1_addr[1]&r_0_addr[12],
r_2_addr[6]&r_1_addr[1]&r_0_addr[11],
r_2_addr[6]&r_1_addr[1]&r_0_addr[10],
r_2_addr[6]&r_1_addr[1]&r_0_addr[9],
r_2_addr[6]&r_1_addr[1]&r_0_addr[8],
r_2_addr[6]&r_1_addr[1]&r_0_addr[7],
r_2_addr[6]&r_1_addr[1]&r_0_addr[6],
r_2_addr[6]&r_1_addr[1]&r_0_addr[5],
r_2_addr[6]&r_1_addr[1]&r_0_addr[4],
r_2_addr[6]&r_1_addr[1]&r_0_addr[3],
r_2_addr[6]&r_1_addr[1]&r_0_addr[2],
r_2_addr[6]&r_1_addr[1]&r_0_addr[1],
r_2_addr[6]&r_1_addr[1]&r_0_addr[0],
r_2_addr[6]&r_1_addr[0]&r_0_addr[15],
r_2_addr[6]&r_1_addr[0]&r_0_addr[14],
r_2_addr[6]&r_1_addr[0]&r_0_addr[13],
r_2_addr[6]&r_1_addr[0]&r_0_addr[12],
r_2_addr[6]&r_1_addr[0]&r_0_addr[11],
r_2_addr[6]&r_1_addr[0]&r_0_addr[10],
r_2_addr[6]&r_1_addr[0]&r_0_addr[9],
r_2_addr[6]&r_1_addr[0]&r_0_addr[8],
r_2_addr[6]&r_1_addr[0]&r_0_addr[7],
r_2_addr[6]&r_1_addr[0]&r_0_addr[6],
r_2_addr[6]&r_1_addr[0]&r_0_addr[5],
r_2_addr[6]&r_1_addr[0]&r_0_addr[4],
r_2_addr[6]&r_1_addr[0]&r_0_addr[3],
r_2_addr[6]&r_1_addr[0]&r_0_addr[2],
r_2_addr[6]&r_1_addr[0]&r_0_addr[1],
r_2_addr[6]&r_1_addr[0]&r_0_addr[0],
r_2_addr[5]&r_1_addr[15]&r_0_addr[15],
r_2_addr[5]&r_1_addr[15]&r_0_addr[14],
r_2_addr[5]&r_1_addr[15]&r_0_addr[13],
r_2_addr[5]&r_1_addr[15]&r_0_addr[12],
r_2_addr[5]&r_1_addr[15]&r_0_addr[11],
r_2_addr[5]&r_1_addr[15]&r_0_addr[10],
r_2_addr[5]&r_1_addr[15]&r_0_addr[9],
r_2_addr[5]&r_1_addr[15]&r_0_addr[8],
r_2_addr[5]&r_1_addr[15]&r_0_addr[7],
r_2_addr[5]&r_1_addr[15]&r_0_addr[6],
r_2_addr[5]&r_1_addr[15]&r_0_addr[5],
r_2_addr[5]&r_1_addr[15]&r_0_addr[4],
r_2_addr[5]&r_1_addr[15]&r_0_addr[3],
r_2_addr[5]&r_1_addr[15]&r_0_addr[2],
r_2_addr[5]&r_1_addr[15]&r_0_addr[1],
r_2_addr[5]&r_1_addr[15]&r_0_addr[0],
r_2_addr[5]&r_1_addr[14]&r_0_addr[15],
r_2_addr[5]&r_1_addr[14]&r_0_addr[14],
r_2_addr[5]&r_1_addr[14]&r_0_addr[13],
r_2_addr[5]&r_1_addr[14]&r_0_addr[12],
r_2_addr[5]&r_1_addr[14]&r_0_addr[11],
r_2_addr[5]&r_1_addr[14]&r_0_addr[10],
r_2_addr[5]&r_1_addr[14]&r_0_addr[9],
r_2_addr[5]&r_1_addr[14]&r_0_addr[8],
r_2_addr[5]&r_1_addr[14]&r_0_addr[7],
r_2_addr[5]&r_1_addr[14]&r_0_addr[6],
r_2_addr[5]&r_1_addr[14]&r_0_addr[5],
r_2_addr[5]&r_1_addr[14]&r_0_addr[4],
r_2_addr[5]&r_1_addr[14]&r_0_addr[3],
r_2_addr[5]&r_1_addr[14]&r_0_addr[2],
r_2_addr[5]&r_1_addr[14]&r_0_addr[1],
r_2_addr[5]&r_1_addr[14]&r_0_addr[0],
r_2_addr[5]&r_1_addr[13]&r_0_addr[15],
r_2_addr[5]&r_1_addr[13]&r_0_addr[14],
r_2_addr[5]&r_1_addr[13]&r_0_addr[13],
r_2_addr[5]&r_1_addr[13]&r_0_addr[12],
r_2_addr[5]&r_1_addr[13]&r_0_addr[11],
r_2_addr[5]&r_1_addr[13]&r_0_addr[10],
r_2_addr[5]&r_1_addr[13]&r_0_addr[9],
r_2_addr[5]&r_1_addr[13]&r_0_addr[8],
r_2_addr[5]&r_1_addr[13]&r_0_addr[7],
r_2_addr[5]&r_1_addr[13]&r_0_addr[6],
r_2_addr[5]&r_1_addr[13]&r_0_addr[5],
r_2_addr[5]&r_1_addr[13]&r_0_addr[4],
r_2_addr[5]&r_1_addr[13]&r_0_addr[3],
r_2_addr[5]&r_1_addr[13]&r_0_addr[2],
r_2_addr[5]&r_1_addr[13]&r_0_addr[1],
r_2_addr[5]&r_1_addr[13]&r_0_addr[0],
r_2_addr[5]&r_1_addr[12]&r_0_addr[15],
r_2_addr[5]&r_1_addr[12]&r_0_addr[14],
r_2_addr[5]&r_1_addr[12]&r_0_addr[13],
r_2_addr[5]&r_1_addr[12]&r_0_addr[12],
r_2_addr[5]&r_1_addr[12]&r_0_addr[11],
r_2_addr[5]&r_1_addr[12]&r_0_addr[10],
r_2_addr[5]&r_1_addr[12]&r_0_addr[9],
r_2_addr[5]&r_1_addr[12]&r_0_addr[8],
r_2_addr[5]&r_1_addr[12]&r_0_addr[7],
r_2_addr[5]&r_1_addr[12]&r_0_addr[6],
r_2_addr[5]&r_1_addr[12]&r_0_addr[5],
r_2_addr[5]&r_1_addr[12]&r_0_addr[4],
r_2_addr[5]&r_1_addr[12]&r_0_addr[3],
r_2_addr[5]&r_1_addr[12]&r_0_addr[2],
r_2_addr[5]&r_1_addr[12]&r_0_addr[1],
r_2_addr[5]&r_1_addr[12]&r_0_addr[0],
r_2_addr[5]&r_1_addr[11]&r_0_addr[15],
r_2_addr[5]&r_1_addr[11]&r_0_addr[14],
r_2_addr[5]&r_1_addr[11]&r_0_addr[13],
r_2_addr[5]&r_1_addr[11]&r_0_addr[12],
r_2_addr[5]&r_1_addr[11]&r_0_addr[11],
r_2_addr[5]&r_1_addr[11]&r_0_addr[10],
r_2_addr[5]&r_1_addr[11]&r_0_addr[9],
r_2_addr[5]&r_1_addr[11]&r_0_addr[8],
r_2_addr[5]&r_1_addr[11]&r_0_addr[7],
r_2_addr[5]&r_1_addr[11]&r_0_addr[6],
r_2_addr[5]&r_1_addr[11]&r_0_addr[5],
r_2_addr[5]&r_1_addr[11]&r_0_addr[4],
r_2_addr[5]&r_1_addr[11]&r_0_addr[3],
r_2_addr[5]&r_1_addr[11]&r_0_addr[2],
r_2_addr[5]&r_1_addr[11]&r_0_addr[1],
r_2_addr[5]&r_1_addr[11]&r_0_addr[0],
r_2_addr[5]&r_1_addr[10]&r_0_addr[15],
r_2_addr[5]&r_1_addr[10]&r_0_addr[14],
r_2_addr[5]&r_1_addr[10]&r_0_addr[13],
r_2_addr[5]&r_1_addr[10]&r_0_addr[12],
r_2_addr[5]&r_1_addr[10]&r_0_addr[11],
r_2_addr[5]&r_1_addr[10]&r_0_addr[10],
r_2_addr[5]&r_1_addr[10]&r_0_addr[9],
r_2_addr[5]&r_1_addr[10]&r_0_addr[8],
r_2_addr[5]&r_1_addr[10]&r_0_addr[7],
r_2_addr[5]&r_1_addr[10]&r_0_addr[6],
r_2_addr[5]&r_1_addr[10]&r_0_addr[5],
r_2_addr[5]&r_1_addr[10]&r_0_addr[4],
r_2_addr[5]&r_1_addr[10]&r_0_addr[3],
r_2_addr[5]&r_1_addr[10]&r_0_addr[2],
r_2_addr[5]&r_1_addr[10]&r_0_addr[1],
r_2_addr[5]&r_1_addr[10]&r_0_addr[0],
r_2_addr[5]&r_1_addr[9]&r_0_addr[15],
r_2_addr[5]&r_1_addr[9]&r_0_addr[14],
r_2_addr[5]&r_1_addr[9]&r_0_addr[13],
r_2_addr[5]&r_1_addr[9]&r_0_addr[12],
r_2_addr[5]&r_1_addr[9]&r_0_addr[11],
r_2_addr[5]&r_1_addr[9]&r_0_addr[10],
r_2_addr[5]&r_1_addr[9]&r_0_addr[9],
r_2_addr[5]&r_1_addr[9]&r_0_addr[8],
r_2_addr[5]&r_1_addr[9]&r_0_addr[7],
r_2_addr[5]&r_1_addr[9]&r_0_addr[6],
r_2_addr[5]&r_1_addr[9]&r_0_addr[5],
r_2_addr[5]&r_1_addr[9]&r_0_addr[4],
r_2_addr[5]&r_1_addr[9]&r_0_addr[3],
r_2_addr[5]&r_1_addr[9]&r_0_addr[2],
r_2_addr[5]&r_1_addr[9]&r_0_addr[1],
r_2_addr[5]&r_1_addr[9]&r_0_addr[0],
r_2_addr[5]&r_1_addr[8]&r_0_addr[15],
r_2_addr[5]&r_1_addr[8]&r_0_addr[14],
r_2_addr[5]&r_1_addr[8]&r_0_addr[13],
r_2_addr[5]&r_1_addr[8]&r_0_addr[12],
r_2_addr[5]&r_1_addr[8]&r_0_addr[11],
r_2_addr[5]&r_1_addr[8]&r_0_addr[10],
r_2_addr[5]&r_1_addr[8]&r_0_addr[9],
r_2_addr[5]&r_1_addr[8]&r_0_addr[8],
r_2_addr[5]&r_1_addr[8]&r_0_addr[7],
r_2_addr[5]&r_1_addr[8]&r_0_addr[6],
r_2_addr[5]&r_1_addr[8]&r_0_addr[5],
r_2_addr[5]&r_1_addr[8]&r_0_addr[4],
r_2_addr[5]&r_1_addr[8]&r_0_addr[3],
r_2_addr[5]&r_1_addr[8]&r_0_addr[2],
r_2_addr[5]&r_1_addr[8]&r_0_addr[1],
r_2_addr[5]&r_1_addr[8]&r_0_addr[0],
r_2_addr[5]&r_1_addr[7]&r_0_addr[15],
r_2_addr[5]&r_1_addr[7]&r_0_addr[14],
r_2_addr[5]&r_1_addr[7]&r_0_addr[13],
r_2_addr[5]&r_1_addr[7]&r_0_addr[12],
r_2_addr[5]&r_1_addr[7]&r_0_addr[11],
r_2_addr[5]&r_1_addr[7]&r_0_addr[10],
r_2_addr[5]&r_1_addr[7]&r_0_addr[9],
r_2_addr[5]&r_1_addr[7]&r_0_addr[8],
r_2_addr[5]&r_1_addr[7]&r_0_addr[7],
r_2_addr[5]&r_1_addr[7]&r_0_addr[6],
r_2_addr[5]&r_1_addr[7]&r_0_addr[5],
r_2_addr[5]&r_1_addr[7]&r_0_addr[4],
r_2_addr[5]&r_1_addr[7]&r_0_addr[3],
r_2_addr[5]&r_1_addr[7]&r_0_addr[2],
r_2_addr[5]&r_1_addr[7]&r_0_addr[1],
r_2_addr[5]&r_1_addr[7]&r_0_addr[0],
r_2_addr[5]&r_1_addr[6]&r_0_addr[15],
r_2_addr[5]&r_1_addr[6]&r_0_addr[14],
r_2_addr[5]&r_1_addr[6]&r_0_addr[13],
r_2_addr[5]&r_1_addr[6]&r_0_addr[12],
r_2_addr[5]&r_1_addr[6]&r_0_addr[11],
r_2_addr[5]&r_1_addr[6]&r_0_addr[10],
r_2_addr[5]&r_1_addr[6]&r_0_addr[9],
r_2_addr[5]&r_1_addr[6]&r_0_addr[8],
r_2_addr[5]&r_1_addr[6]&r_0_addr[7],
r_2_addr[5]&r_1_addr[6]&r_0_addr[6],
r_2_addr[5]&r_1_addr[6]&r_0_addr[5],
r_2_addr[5]&r_1_addr[6]&r_0_addr[4],
r_2_addr[5]&r_1_addr[6]&r_0_addr[3],
r_2_addr[5]&r_1_addr[6]&r_0_addr[2],
r_2_addr[5]&r_1_addr[6]&r_0_addr[1],
r_2_addr[5]&r_1_addr[6]&r_0_addr[0],
r_2_addr[5]&r_1_addr[5]&r_0_addr[15],
r_2_addr[5]&r_1_addr[5]&r_0_addr[14],
r_2_addr[5]&r_1_addr[5]&r_0_addr[13],
r_2_addr[5]&r_1_addr[5]&r_0_addr[12],
r_2_addr[5]&r_1_addr[5]&r_0_addr[11],
r_2_addr[5]&r_1_addr[5]&r_0_addr[10],
r_2_addr[5]&r_1_addr[5]&r_0_addr[9],
r_2_addr[5]&r_1_addr[5]&r_0_addr[8],
r_2_addr[5]&r_1_addr[5]&r_0_addr[7],
r_2_addr[5]&r_1_addr[5]&r_0_addr[6],
r_2_addr[5]&r_1_addr[5]&r_0_addr[5],
r_2_addr[5]&r_1_addr[5]&r_0_addr[4],
r_2_addr[5]&r_1_addr[5]&r_0_addr[3],
r_2_addr[5]&r_1_addr[5]&r_0_addr[2],
r_2_addr[5]&r_1_addr[5]&r_0_addr[1],
r_2_addr[5]&r_1_addr[5]&r_0_addr[0],
r_2_addr[5]&r_1_addr[4]&r_0_addr[15],
r_2_addr[5]&r_1_addr[4]&r_0_addr[14],
r_2_addr[5]&r_1_addr[4]&r_0_addr[13],
r_2_addr[5]&r_1_addr[4]&r_0_addr[12],
r_2_addr[5]&r_1_addr[4]&r_0_addr[11],
r_2_addr[5]&r_1_addr[4]&r_0_addr[10],
r_2_addr[5]&r_1_addr[4]&r_0_addr[9],
r_2_addr[5]&r_1_addr[4]&r_0_addr[8],
r_2_addr[5]&r_1_addr[4]&r_0_addr[7],
r_2_addr[5]&r_1_addr[4]&r_0_addr[6],
r_2_addr[5]&r_1_addr[4]&r_0_addr[5],
r_2_addr[5]&r_1_addr[4]&r_0_addr[4],
r_2_addr[5]&r_1_addr[4]&r_0_addr[3],
r_2_addr[5]&r_1_addr[4]&r_0_addr[2],
r_2_addr[5]&r_1_addr[4]&r_0_addr[1],
r_2_addr[5]&r_1_addr[4]&r_0_addr[0],
r_2_addr[5]&r_1_addr[3]&r_0_addr[15],
r_2_addr[5]&r_1_addr[3]&r_0_addr[14],
r_2_addr[5]&r_1_addr[3]&r_0_addr[13],
r_2_addr[5]&r_1_addr[3]&r_0_addr[12],
r_2_addr[5]&r_1_addr[3]&r_0_addr[11],
r_2_addr[5]&r_1_addr[3]&r_0_addr[10],
r_2_addr[5]&r_1_addr[3]&r_0_addr[9],
r_2_addr[5]&r_1_addr[3]&r_0_addr[8],
r_2_addr[5]&r_1_addr[3]&r_0_addr[7],
r_2_addr[5]&r_1_addr[3]&r_0_addr[6],
r_2_addr[5]&r_1_addr[3]&r_0_addr[5],
r_2_addr[5]&r_1_addr[3]&r_0_addr[4],
r_2_addr[5]&r_1_addr[3]&r_0_addr[3],
r_2_addr[5]&r_1_addr[3]&r_0_addr[2],
r_2_addr[5]&r_1_addr[3]&r_0_addr[1],
r_2_addr[5]&r_1_addr[3]&r_0_addr[0],
r_2_addr[5]&r_1_addr[2]&r_0_addr[15],
r_2_addr[5]&r_1_addr[2]&r_0_addr[14],
r_2_addr[5]&r_1_addr[2]&r_0_addr[13],
r_2_addr[5]&r_1_addr[2]&r_0_addr[12],
r_2_addr[5]&r_1_addr[2]&r_0_addr[11],
r_2_addr[5]&r_1_addr[2]&r_0_addr[10],
r_2_addr[5]&r_1_addr[2]&r_0_addr[9],
r_2_addr[5]&r_1_addr[2]&r_0_addr[8],
r_2_addr[5]&r_1_addr[2]&r_0_addr[7],
r_2_addr[5]&r_1_addr[2]&r_0_addr[6],
r_2_addr[5]&r_1_addr[2]&r_0_addr[5],
r_2_addr[5]&r_1_addr[2]&r_0_addr[4],
r_2_addr[5]&r_1_addr[2]&r_0_addr[3],
r_2_addr[5]&r_1_addr[2]&r_0_addr[2],
r_2_addr[5]&r_1_addr[2]&r_0_addr[1],
r_2_addr[5]&r_1_addr[2]&r_0_addr[0],
r_2_addr[5]&r_1_addr[1]&r_0_addr[15],
r_2_addr[5]&r_1_addr[1]&r_0_addr[14],
r_2_addr[5]&r_1_addr[1]&r_0_addr[13],
r_2_addr[5]&r_1_addr[1]&r_0_addr[12],
r_2_addr[5]&r_1_addr[1]&r_0_addr[11],
r_2_addr[5]&r_1_addr[1]&r_0_addr[10],
r_2_addr[5]&r_1_addr[1]&r_0_addr[9],
r_2_addr[5]&r_1_addr[1]&r_0_addr[8],
r_2_addr[5]&r_1_addr[1]&r_0_addr[7],
r_2_addr[5]&r_1_addr[1]&r_0_addr[6],
r_2_addr[5]&r_1_addr[1]&r_0_addr[5],
r_2_addr[5]&r_1_addr[1]&r_0_addr[4],
r_2_addr[5]&r_1_addr[1]&r_0_addr[3],
r_2_addr[5]&r_1_addr[1]&r_0_addr[2],
r_2_addr[5]&r_1_addr[1]&r_0_addr[1],
r_2_addr[5]&r_1_addr[1]&r_0_addr[0],
r_2_addr[5]&r_1_addr[0]&r_0_addr[15],
r_2_addr[5]&r_1_addr[0]&r_0_addr[14],
r_2_addr[5]&r_1_addr[0]&r_0_addr[13],
r_2_addr[5]&r_1_addr[0]&r_0_addr[12],
r_2_addr[5]&r_1_addr[0]&r_0_addr[11],
r_2_addr[5]&r_1_addr[0]&r_0_addr[10],
r_2_addr[5]&r_1_addr[0]&r_0_addr[9],
r_2_addr[5]&r_1_addr[0]&r_0_addr[8],
r_2_addr[5]&r_1_addr[0]&r_0_addr[7],
r_2_addr[5]&r_1_addr[0]&r_0_addr[6],
r_2_addr[5]&r_1_addr[0]&r_0_addr[5],
r_2_addr[5]&r_1_addr[0]&r_0_addr[4],
r_2_addr[5]&r_1_addr[0]&r_0_addr[3],
r_2_addr[5]&r_1_addr[0]&r_0_addr[2],
r_2_addr[5]&r_1_addr[0]&r_0_addr[1],
r_2_addr[5]&r_1_addr[0]&r_0_addr[0],
r_2_addr[4]&r_1_addr[15]&r_0_addr[15],
r_2_addr[4]&r_1_addr[15]&r_0_addr[14],
r_2_addr[4]&r_1_addr[15]&r_0_addr[13],
r_2_addr[4]&r_1_addr[15]&r_0_addr[12],
r_2_addr[4]&r_1_addr[15]&r_0_addr[11],
r_2_addr[4]&r_1_addr[15]&r_0_addr[10],
r_2_addr[4]&r_1_addr[15]&r_0_addr[9],
r_2_addr[4]&r_1_addr[15]&r_0_addr[8],
r_2_addr[4]&r_1_addr[15]&r_0_addr[7],
r_2_addr[4]&r_1_addr[15]&r_0_addr[6],
r_2_addr[4]&r_1_addr[15]&r_0_addr[5],
r_2_addr[4]&r_1_addr[15]&r_0_addr[4],
r_2_addr[4]&r_1_addr[15]&r_0_addr[3],
r_2_addr[4]&r_1_addr[15]&r_0_addr[2],
r_2_addr[4]&r_1_addr[15]&r_0_addr[1],
r_2_addr[4]&r_1_addr[15]&r_0_addr[0],
r_2_addr[4]&r_1_addr[14]&r_0_addr[15],
r_2_addr[4]&r_1_addr[14]&r_0_addr[14],
r_2_addr[4]&r_1_addr[14]&r_0_addr[13],
r_2_addr[4]&r_1_addr[14]&r_0_addr[12],
r_2_addr[4]&r_1_addr[14]&r_0_addr[11],
r_2_addr[4]&r_1_addr[14]&r_0_addr[10],
r_2_addr[4]&r_1_addr[14]&r_0_addr[9],
r_2_addr[4]&r_1_addr[14]&r_0_addr[8],
r_2_addr[4]&r_1_addr[14]&r_0_addr[7],
r_2_addr[4]&r_1_addr[14]&r_0_addr[6],
r_2_addr[4]&r_1_addr[14]&r_0_addr[5],
r_2_addr[4]&r_1_addr[14]&r_0_addr[4],
r_2_addr[4]&r_1_addr[14]&r_0_addr[3],
r_2_addr[4]&r_1_addr[14]&r_0_addr[2],
r_2_addr[4]&r_1_addr[14]&r_0_addr[1],
r_2_addr[4]&r_1_addr[14]&r_0_addr[0],
r_2_addr[4]&r_1_addr[13]&r_0_addr[15],
r_2_addr[4]&r_1_addr[13]&r_0_addr[14],
r_2_addr[4]&r_1_addr[13]&r_0_addr[13],
r_2_addr[4]&r_1_addr[13]&r_0_addr[12],
r_2_addr[4]&r_1_addr[13]&r_0_addr[11],
r_2_addr[4]&r_1_addr[13]&r_0_addr[10],
r_2_addr[4]&r_1_addr[13]&r_0_addr[9],
r_2_addr[4]&r_1_addr[13]&r_0_addr[8],
r_2_addr[4]&r_1_addr[13]&r_0_addr[7],
r_2_addr[4]&r_1_addr[13]&r_0_addr[6],
r_2_addr[4]&r_1_addr[13]&r_0_addr[5],
r_2_addr[4]&r_1_addr[13]&r_0_addr[4],
r_2_addr[4]&r_1_addr[13]&r_0_addr[3],
r_2_addr[4]&r_1_addr[13]&r_0_addr[2],
r_2_addr[4]&r_1_addr[13]&r_0_addr[1],
r_2_addr[4]&r_1_addr[13]&r_0_addr[0],
r_2_addr[4]&r_1_addr[12]&r_0_addr[15],
r_2_addr[4]&r_1_addr[12]&r_0_addr[14],
r_2_addr[4]&r_1_addr[12]&r_0_addr[13],
r_2_addr[4]&r_1_addr[12]&r_0_addr[12],
r_2_addr[4]&r_1_addr[12]&r_0_addr[11],
r_2_addr[4]&r_1_addr[12]&r_0_addr[10],
r_2_addr[4]&r_1_addr[12]&r_0_addr[9],
r_2_addr[4]&r_1_addr[12]&r_0_addr[8],
r_2_addr[4]&r_1_addr[12]&r_0_addr[7],
r_2_addr[4]&r_1_addr[12]&r_0_addr[6],
r_2_addr[4]&r_1_addr[12]&r_0_addr[5],
r_2_addr[4]&r_1_addr[12]&r_0_addr[4],
r_2_addr[4]&r_1_addr[12]&r_0_addr[3],
r_2_addr[4]&r_1_addr[12]&r_0_addr[2],
r_2_addr[4]&r_1_addr[12]&r_0_addr[1],
r_2_addr[4]&r_1_addr[12]&r_0_addr[0],
r_2_addr[4]&r_1_addr[11]&r_0_addr[15],
r_2_addr[4]&r_1_addr[11]&r_0_addr[14],
r_2_addr[4]&r_1_addr[11]&r_0_addr[13],
r_2_addr[4]&r_1_addr[11]&r_0_addr[12],
r_2_addr[4]&r_1_addr[11]&r_0_addr[11],
r_2_addr[4]&r_1_addr[11]&r_0_addr[10],
r_2_addr[4]&r_1_addr[11]&r_0_addr[9],
r_2_addr[4]&r_1_addr[11]&r_0_addr[8],
r_2_addr[4]&r_1_addr[11]&r_0_addr[7],
r_2_addr[4]&r_1_addr[11]&r_0_addr[6],
r_2_addr[4]&r_1_addr[11]&r_0_addr[5],
r_2_addr[4]&r_1_addr[11]&r_0_addr[4],
r_2_addr[4]&r_1_addr[11]&r_0_addr[3],
r_2_addr[4]&r_1_addr[11]&r_0_addr[2],
r_2_addr[4]&r_1_addr[11]&r_0_addr[1],
r_2_addr[4]&r_1_addr[11]&r_0_addr[0],
r_2_addr[4]&r_1_addr[10]&r_0_addr[15],
r_2_addr[4]&r_1_addr[10]&r_0_addr[14],
r_2_addr[4]&r_1_addr[10]&r_0_addr[13],
r_2_addr[4]&r_1_addr[10]&r_0_addr[12],
r_2_addr[4]&r_1_addr[10]&r_0_addr[11],
r_2_addr[4]&r_1_addr[10]&r_0_addr[10],
r_2_addr[4]&r_1_addr[10]&r_0_addr[9],
r_2_addr[4]&r_1_addr[10]&r_0_addr[8],
r_2_addr[4]&r_1_addr[10]&r_0_addr[7],
r_2_addr[4]&r_1_addr[10]&r_0_addr[6],
r_2_addr[4]&r_1_addr[10]&r_0_addr[5],
r_2_addr[4]&r_1_addr[10]&r_0_addr[4],
r_2_addr[4]&r_1_addr[10]&r_0_addr[3],
r_2_addr[4]&r_1_addr[10]&r_0_addr[2],
r_2_addr[4]&r_1_addr[10]&r_0_addr[1],
r_2_addr[4]&r_1_addr[10]&r_0_addr[0],
r_2_addr[4]&r_1_addr[9]&r_0_addr[15],
r_2_addr[4]&r_1_addr[9]&r_0_addr[14],
r_2_addr[4]&r_1_addr[9]&r_0_addr[13],
r_2_addr[4]&r_1_addr[9]&r_0_addr[12],
r_2_addr[4]&r_1_addr[9]&r_0_addr[11],
r_2_addr[4]&r_1_addr[9]&r_0_addr[10],
r_2_addr[4]&r_1_addr[9]&r_0_addr[9],
r_2_addr[4]&r_1_addr[9]&r_0_addr[8],
r_2_addr[4]&r_1_addr[9]&r_0_addr[7],
r_2_addr[4]&r_1_addr[9]&r_0_addr[6],
r_2_addr[4]&r_1_addr[9]&r_0_addr[5],
r_2_addr[4]&r_1_addr[9]&r_0_addr[4],
r_2_addr[4]&r_1_addr[9]&r_0_addr[3],
r_2_addr[4]&r_1_addr[9]&r_0_addr[2],
r_2_addr[4]&r_1_addr[9]&r_0_addr[1],
r_2_addr[4]&r_1_addr[9]&r_0_addr[0],
r_2_addr[4]&r_1_addr[8]&r_0_addr[15],
r_2_addr[4]&r_1_addr[8]&r_0_addr[14],
r_2_addr[4]&r_1_addr[8]&r_0_addr[13],
r_2_addr[4]&r_1_addr[8]&r_0_addr[12],
r_2_addr[4]&r_1_addr[8]&r_0_addr[11],
r_2_addr[4]&r_1_addr[8]&r_0_addr[10],
r_2_addr[4]&r_1_addr[8]&r_0_addr[9],
r_2_addr[4]&r_1_addr[8]&r_0_addr[8],
r_2_addr[4]&r_1_addr[8]&r_0_addr[7],
r_2_addr[4]&r_1_addr[8]&r_0_addr[6],
r_2_addr[4]&r_1_addr[8]&r_0_addr[5],
r_2_addr[4]&r_1_addr[8]&r_0_addr[4],
r_2_addr[4]&r_1_addr[8]&r_0_addr[3],
r_2_addr[4]&r_1_addr[8]&r_0_addr[2],
r_2_addr[4]&r_1_addr[8]&r_0_addr[1],
r_2_addr[4]&r_1_addr[8]&r_0_addr[0],
r_2_addr[4]&r_1_addr[7]&r_0_addr[15],
r_2_addr[4]&r_1_addr[7]&r_0_addr[14],
r_2_addr[4]&r_1_addr[7]&r_0_addr[13],
r_2_addr[4]&r_1_addr[7]&r_0_addr[12],
r_2_addr[4]&r_1_addr[7]&r_0_addr[11],
r_2_addr[4]&r_1_addr[7]&r_0_addr[10],
r_2_addr[4]&r_1_addr[7]&r_0_addr[9],
r_2_addr[4]&r_1_addr[7]&r_0_addr[8],
r_2_addr[4]&r_1_addr[7]&r_0_addr[7],
r_2_addr[4]&r_1_addr[7]&r_0_addr[6],
r_2_addr[4]&r_1_addr[7]&r_0_addr[5],
r_2_addr[4]&r_1_addr[7]&r_0_addr[4],
r_2_addr[4]&r_1_addr[7]&r_0_addr[3],
r_2_addr[4]&r_1_addr[7]&r_0_addr[2],
r_2_addr[4]&r_1_addr[7]&r_0_addr[1],
r_2_addr[4]&r_1_addr[7]&r_0_addr[0],
r_2_addr[4]&r_1_addr[6]&r_0_addr[15],
r_2_addr[4]&r_1_addr[6]&r_0_addr[14],
r_2_addr[4]&r_1_addr[6]&r_0_addr[13],
r_2_addr[4]&r_1_addr[6]&r_0_addr[12],
r_2_addr[4]&r_1_addr[6]&r_0_addr[11],
r_2_addr[4]&r_1_addr[6]&r_0_addr[10],
r_2_addr[4]&r_1_addr[6]&r_0_addr[9],
r_2_addr[4]&r_1_addr[6]&r_0_addr[8],
r_2_addr[4]&r_1_addr[6]&r_0_addr[7],
r_2_addr[4]&r_1_addr[6]&r_0_addr[6],
r_2_addr[4]&r_1_addr[6]&r_0_addr[5],
r_2_addr[4]&r_1_addr[6]&r_0_addr[4],
r_2_addr[4]&r_1_addr[6]&r_0_addr[3],
r_2_addr[4]&r_1_addr[6]&r_0_addr[2],
r_2_addr[4]&r_1_addr[6]&r_0_addr[1],
r_2_addr[4]&r_1_addr[6]&r_0_addr[0],
r_2_addr[4]&r_1_addr[5]&r_0_addr[15],
r_2_addr[4]&r_1_addr[5]&r_0_addr[14],
r_2_addr[4]&r_1_addr[5]&r_0_addr[13],
r_2_addr[4]&r_1_addr[5]&r_0_addr[12],
r_2_addr[4]&r_1_addr[5]&r_0_addr[11],
r_2_addr[4]&r_1_addr[5]&r_0_addr[10],
r_2_addr[4]&r_1_addr[5]&r_0_addr[9],
r_2_addr[4]&r_1_addr[5]&r_0_addr[8],
r_2_addr[4]&r_1_addr[5]&r_0_addr[7],
r_2_addr[4]&r_1_addr[5]&r_0_addr[6],
r_2_addr[4]&r_1_addr[5]&r_0_addr[5],
r_2_addr[4]&r_1_addr[5]&r_0_addr[4],
r_2_addr[4]&r_1_addr[5]&r_0_addr[3],
r_2_addr[4]&r_1_addr[5]&r_0_addr[2],
r_2_addr[4]&r_1_addr[5]&r_0_addr[1],
r_2_addr[4]&r_1_addr[5]&r_0_addr[0],
r_2_addr[4]&r_1_addr[4]&r_0_addr[15],
r_2_addr[4]&r_1_addr[4]&r_0_addr[14],
r_2_addr[4]&r_1_addr[4]&r_0_addr[13],
r_2_addr[4]&r_1_addr[4]&r_0_addr[12],
r_2_addr[4]&r_1_addr[4]&r_0_addr[11],
r_2_addr[4]&r_1_addr[4]&r_0_addr[10],
r_2_addr[4]&r_1_addr[4]&r_0_addr[9],
r_2_addr[4]&r_1_addr[4]&r_0_addr[8],
r_2_addr[4]&r_1_addr[4]&r_0_addr[7],
r_2_addr[4]&r_1_addr[4]&r_0_addr[6],
r_2_addr[4]&r_1_addr[4]&r_0_addr[5],
r_2_addr[4]&r_1_addr[4]&r_0_addr[4],
r_2_addr[4]&r_1_addr[4]&r_0_addr[3],
r_2_addr[4]&r_1_addr[4]&r_0_addr[2],
r_2_addr[4]&r_1_addr[4]&r_0_addr[1],
r_2_addr[4]&r_1_addr[4]&r_0_addr[0],
r_2_addr[4]&r_1_addr[3]&r_0_addr[15],
r_2_addr[4]&r_1_addr[3]&r_0_addr[14],
r_2_addr[4]&r_1_addr[3]&r_0_addr[13],
r_2_addr[4]&r_1_addr[3]&r_0_addr[12],
r_2_addr[4]&r_1_addr[3]&r_0_addr[11],
r_2_addr[4]&r_1_addr[3]&r_0_addr[10],
r_2_addr[4]&r_1_addr[3]&r_0_addr[9],
r_2_addr[4]&r_1_addr[3]&r_0_addr[8],
r_2_addr[4]&r_1_addr[3]&r_0_addr[7],
r_2_addr[4]&r_1_addr[3]&r_0_addr[6],
r_2_addr[4]&r_1_addr[3]&r_0_addr[5],
r_2_addr[4]&r_1_addr[3]&r_0_addr[4],
r_2_addr[4]&r_1_addr[3]&r_0_addr[3],
r_2_addr[4]&r_1_addr[3]&r_0_addr[2],
r_2_addr[4]&r_1_addr[3]&r_0_addr[1],
r_2_addr[4]&r_1_addr[3]&r_0_addr[0],
r_2_addr[4]&r_1_addr[2]&r_0_addr[15],
r_2_addr[4]&r_1_addr[2]&r_0_addr[14],
r_2_addr[4]&r_1_addr[2]&r_0_addr[13],
r_2_addr[4]&r_1_addr[2]&r_0_addr[12],
r_2_addr[4]&r_1_addr[2]&r_0_addr[11],
r_2_addr[4]&r_1_addr[2]&r_0_addr[10],
r_2_addr[4]&r_1_addr[2]&r_0_addr[9],
r_2_addr[4]&r_1_addr[2]&r_0_addr[8],
r_2_addr[4]&r_1_addr[2]&r_0_addr[7],
r_2_addr[4]&r_1_addr[2]&r_0_addr[6],
r_2_addr[4]&r_1_addr[2]&r_0_addr[5],
r_2_addr[4]&r_1_addr[2]&r_0_addr[4],
r_2_addr[4]&r_1_addr[2]&r_0_addr[3],
r_2_addr[4]&r_1_addr[2]&r_0_addr[2],
r_2_addr[4]&r_1_addr[2]&r_0_addr[1],
r_2_addr[4]&r_1_addr[2]&r_0_addr[0],
r_2_addr[4]&r_1_addr[1]&r_0_addr[15],
r_2_addr[4]&r_1_addr[1]&r_0_addr[14],
r_2_addr[4]&r_1_addr[1]&r_0_addr[13],
r_2_addr[4]&r_1_addr[1]&r_0_addr[12],
r_2_addr[4]&r_1_addr[1]&r_0_addr[11],
r_2_addr[4]&r_1_addr[1]&r_0_addr[10],
r_2_addr[4]&r_1_addr[1]&r_0_addr[9],
r_2_addr[4]&r_1_addr[1]&r_0_addr[8],
r_2_addr[4]&r_1_addr[1]&r_0_addr[7],
r_2_addr[4]&r_1_addr[1]&r_0_addr[6],
r_2_addr[4]&r_1_addr[1]&r_0_addr[5],
r_2_addr[4]&r_1_addr[1]&r_0_addr[4],
r_2_addr[4]&r_1_addr[1]&r_0_addr[3],
r_2_addr[4]&r_1_addr[1]&r_0_addr[2],
r_2_addr[4]&r_1_addr[1]&r_0_addr[1],
r_2_addr[4]&r_1_addr[1]&r_0_addr[0],
r_2_addr[4]&r_1_addr[0]&r_0_addr[15],
r_2_addr[4]&r_1_addr[0]&r_0_addr[14],
r_2_addr[4]&r_1_addr[0]&r_0_addr[13],
r_2_addr[4]&r_1_addr[0]&r_0_addr[12],
r_2_addr[4]&r_1_addr[0]&r_0_addr[11],
r_2_addr[4]&r_1_addr[0]&r_0_addr[10],
r_2_addr[4]&r_1_addr[0]&r_0_addr[9],
r_2_addr[4]&r_1_addr[0]&r_0_addr[8],
r_2_addr[4]&r_1_addr[0]&r_0_addr[7],
r_2_addr[4]&r_1_addr[0]&r_0_addr[6],
r_2_addr[4]&r_1_addr[0]&r_0_addr[5],
r_2_addr[4]&r_1_addr[0]&r_0_addr[4],
r_2_addr[4]&r_1_addr[0]&r_0_addr[3],
r_2_addr[4]&r_1_addr[0]&r_0_addr[2],
r_2_addr[4]&r_1_addr[0]&r_0_addr[1],
r_2_addr[4]&r_1_addr[0]&r_0_addr[0],
r_2_addr[3]&r_1_addr[15]&r_0_addr[15],
r_2_addr[3]&r_1_addr[15]&r_0_addr[14],
r_2_addr[3]&r_1_addr[15]&r_0_addr[13],
r_2_addr[3]&r_1_addr[15]&r_0_addr[12],
r_2_addr[3]&r_1_addr[15]&r_0_addr[11],
r_2_addr[3]&r_1_addr[15]&r_0_addr[10],
r_2_addr[3]&r_1_addr[15]&r_0_addr[9],
r_2_addr[3]&r_1_addr[15]&r_0_addr[8],
r_2_addr[3]&r_1_addr[15]&r_0_addr[7],
r_2_addr[3]&r_1_addr[15]&r_0_addr[6],
r_2_addr[3]&r_1_addr[15]&r_0_addr[5],
r_2_addr[3]&r_1_addr[15]&r_0_addr[4],
r_2_addr[3]&r_1_addr[15]&r_0_addr[3],
r_2_addr[3]&r_1_addr[15]&r_0_addr[2],
r_2_addr[3]&r_1_addr[15]&r_0_addr[1],
r_2_addr[3]&r_1_addr[15]&r_0_addr[0],
r_2_addr[3]&r_1_addr[14]&r_0_addr[15],
r_2_addr[3]&r_1_addr[14]&r_0_addr[14],
r_2_addr[3]&r_1_addr[14]&r_0_addr[13],
r_2_addr[3]&r_1_addr[14]&r_0_addr[12],
r_2_addr[3]&r_1_addr[14]&r_0_addr[11],
r_2_addr[3]&r_1_addr[14]&r_0_addr[10],
r_2_addr[3]&r_1_addr[14]&r_0_addr[9],
r_2_addr[3]&r_1_addr[14]&r_0_addr[8],
r_2_addr[3]&r_1_addr[14]&r_0_addr[7],
r_2_addr[3]&r_1_addr[14]&r_0_addr[6],
r_2_addr[3]&r_1_addr[14]&r_0_addr[5],
r_2_addr[3]&r_1_addr[14]&r_0_addr[4],
r_2_addr[3]&r_1_addr[14]&r_0_addr[3],
r_2_addr[3]&r_1_addr[14]&r_0_addr[2],
r_2_addr[3]&r_1_addr[14]&r_0_addr[1],
r_2_addr[3]&r_1_addr[14]&r_0_addr[0],
r_2_addr[3]&r_1_addr[13]&r_0_addr[15],
r_2_addr[3]&r_1_addr[13]&r_0_addr[14],
r_2_addr[3]&r_1_addr[13]&r_0_addr[13],
r_2_addr[3]&r_1_addr[13]&r_0_addr[12],
r_2_addr[3]&r_1_addr[13]&r_0_addr[11],
r_2_addr[3]&r_1_addr[13]&r_0_addr[10],
r_2_addr[3]&r_1_addr[13]&r_0_addr[9],
r_2_addr[3]&r_1_addr[13]&r_0_addr[8],
r_2_addr[3]&r_1_addr[13]&r_0_addr[7],
r_2_addr[3]&r_1_addr[13]&r_0_addr[6],
r_2_addr[3]&r_1_addr[13]&r_0_addr[5],
r_2_addr[3]&r_1_addr[13]&r_0_addr[4],
r_2_addr[3]&r_1_addr[13]&r_0_addr[3],
r_2_addr[3]&r_1_addr[13]&r_0_addr[2],
r_2_addr[3]&r_1_addr[13]&r_0_addr[1],
r_2_addr[3]&r_1_addr[13]&r_0_addr[0],
r_2_addr[3]&r_1_addr[12]&r_0_addr[15],
r_2_addr[3]&r_1_addr[12]&r_0_addr[14],
r_2_addr[3]&r_1_addr[12]&r_0_addr[13],
r_2_addr[3]&r_1_addr[12]&r_0_addr[12],
r_2_addr[3]&r_1_addr[12]&r_0_addr[11],
r_2_addr[3]&r_1_addr[12]&r_0_addr[10],
r_2_addr[3]&r_1_addr[12]&r_0_addr[9],
r_2_addr[3]&r_1_addr[12]&r_0_addr[8],
r_2_addr[3]&r_1_addr[12]&r_0_addr[7],
r_2_addr[3]&r_1_addr[12]&r_0_addr[6],
r_2_addr[3]&r_1_addr[12]&r_0_addr[5],
r_2_addr[3]&r_1_addr[12]&r_0_addr[4],
r_2_addr[3]&r_1_addr[12]&r_0_addr[3],
r_2_addr[3]&r_1_addr[12]&r_0_addr[2],
r_2_addr[3]&r_1_addr[12]&r_0_addr[1],
r_2_addr[3]&r_1_addr[12]&r_0_addr[0],
r_2_addr[3]&r_1_addr[11]&r_0_addr[15],
r_2_addr[3]&r_1_addr[11]&r_0_addr[14],
r_2_addr[3]&r_1_addr[11]&r_0_addr[13],
r_2_addr[3]&r_1_addr[11]&r_0_addr[12],
r_2_addr[3]&r_1_addr[11]&r_0_addr[11],
r_2_addr[3]&r_1_addr[11]&r_0_addr[10],
r_2_addr[3]&r_1_addr[11]&r_0_addr[9],
r_2_addr[3]&r_1_addr[11]&r_0_addr[8],
r_2_addr[3]&r_1_addr[11]&r_0_addr[7],
r_2_addr[3]&r_1_addr[11]&r_0_addr[6],
r_2_addr[3]&r_1_addr[11]&r_0_addr[5],
r_2_addr[3]&r_1_addr[11]&r_0_addr[4],
r_2_addr[3]&r_1_addr[11]&r_0_addr[3],
r_2_addr[3]&r_1_addr[11]&r_0_addr[2],
r_2_addr[3]&r_1_addr[11]&r_0_addr[1],
r_2_addr[3]&r_1_addr[11]&r_0_addr[0],
r_2_addr[3]&r_1_addr[10]&r_0_addr[15],
r_2_addr[3]&r_1_addr[10]&r_0_addr[14],
r_2_addr[3]&r_1_addr[10]&r_0_addr[13],
r_2_addr[3]&r_1_addr[10]&r_0_addr[12],
r_2_addr[3]&r_1_addr[10]&r_0_addr[11],
r_2_addr[3]&r_1_addr[10]&r_0_addr[10],
r_2_addr[3]&r_1_addr[10]&r_0_addr[9],
r_2_addr[3]&r_1_addr[10]&r_0_addr[8],
r_2_addr[3]&r_1_addr[10]&r_0_addr[7],
r_2_addr[3]&r_1_addr[10]&r_0_addr[6],
r_2_addr[3]&r_1_addr[10]&r_0_addr[5],
r_2_addr[3]&r_1_addr[10]&r_0_addr[4],
r_2_addr[3]&r_1_addr[10]&r_0_addr[3],
r_2_addr[3]&r_1_addr[10]&r_0_addr[2],
r_2_addr[3]&r_1_addr[10]&r_0_addr[1],
r_2_addr[3]&r_1_addr[10]&r_0_addr[0],
r_2_addr[3]&r_1_addr[9]&r_0_addr[15],
r_2_addr[3]&r_1_addr[9]&r_0_addr[14],
r_2_addr[3]&r_1_addr[9]&r_0_addr[13],
r_2_addr[3]&r_1_addr[9]&r_0_addr[12],
r_2_addr[3]&r_1_addr[9]&r_0_addr[11],
r_2_addr[3]&r_1_addr[9]&r_0_addr[10],
r_2_addr[3]&r_1_addr[9]&r_0_addr[9],
r_2_addr[3]&r_1_addr[9]&r_0_addr[8],
r_2_addr[3]&r_1_addr[9]&r_0_addr[7],
r_2_addr[3]&r_1_addr[9]&r_0_addr[6],
r_2_addr[3]&r_1_addr[9]&r_0_addr[5],
r_2_addr[3]&r_1_addr[9]&r_0_addr[4],
r_2_addr[3]&r_1_addr[9]&r_0_addr[3],
r_2_addr[3]&r_1_addr[9]&r_0_addr[2],
r_2_addr[3]&r_1_addr[9]&r_0_addr[1],
r_2_addr[3]&r_1_addr[9]&r_0_addr[0],
r_2_addr[3]&r_1_addr[8]&r_0_addr[15],
r_2_addr[3]&r_1_addr[8]&r_0_addr[14],
r_2_addr[3]&r_1_addr[8]&r_0_addr[13],
r_2_addr[3]&r_1_addr[8]&r_0_addr[12],
r_2_addr[3]&r_1_addr[8]&r_0_addr[11],
r_2_addr[3]&r_1_addr[8]&r_0_addr[10],
r_2_addr[3]&r_1_addr[8]&r_0_addr[9],
r_2_addr[3]&r_1_addr[8]&r_0_addr[8],
r_2_addr[3]&r_1_addr[8]&r_0_addr[7],
r_2_addr[3]&r_1_addr[8]&r_0_addr[6],
r_2_addr[3]&r_1_addr[8]&r_0_addr[5],
r_2_addr[3]&r_1_addr[8]&r_0_addr[4],
r_2_addr[3]&r_1_addr[8]&r_0_addr[3],
r_2_addr[3]&r_1_addr[8]&r_0_addr[2],
r_2_addr[3]&r_1_addr[8]&r_0_addr[1],
r_2_addr[3]&r_1_addr[8]&r_0_addr[0],
r_2_addr[3]&r_1_addr[7]&r_0_addr[15],
r_2_addr[3]&r_1_addr[7]&r_0_addr[14],
r_2_addr[3]&r_1_addr[7]&r_0_addr[13],
r_2_addr[3]&r_1_addr[7]&r_0_addr[12],
r_2_addr[3]&r_1_addr[7]&r_0_addr[11],
r_2_addr[3]&r_1_addr[7]&r_0_addr[10],
r_2_addr[3]&r_1_addr[7]&r_0_addr[9],
r_2_addr[3]&r_1_addr[7]&r_0_addr[8],
r_2_addr[3]&r_1_addr[7]&r_0_addr[7],
r_2_addr[3]&r_1_addr[7]&r_0_addr[6],
r_2_addr[3]&r_1_addr[7]&r_0_addr[5],
r_2_addr[3]&r_1_addr[7]&r_0_addr[4],
r_2_addr[3]&r_1_addr[7]&r_0_addr[3],
r_2_addr[3]&r_1_addr[7]&r_0_addr[2],
r_2_addr[3]&r_1_addr[7]&r_0_addr[1],
r_2_addr[3]&r_1_addr[7]&r_0_addr[0],
r_2_addr[3]&r_1_addr[6]&r_0_addr[15],
r_2_addr[3]&r_1_addr[6]&r_0_addr[14],
r_2_addr[3]&r_1_addr[6]&r_0_addr[13],
r_2_addr[3]&r_1_addr[6]&r_0_addr[12],
r_2_addr[3]&r_1_addr[6]&r_0_addr[11],
r_2_addr[3]&r_1_addr[6]&r_0_addr[10],
r_2_addr[3]&r_1_addr[6]&r_0_addr[9],
r_2_addr[3]&r_1_addr[6]&r_0_addr[8],
r_2_addr[3]&r_1_addr[6]&r_0_addr[7],
r_2_addr[3]&r_1_addr[6]&r_0_addr[6],
r_2_addr[3]&r_1_addr[6]&r_0_addr[5],
r_2_addr[3]&r_1_addr[6]&r_0_addr[4],
r_2_addr[3]&r_1_addr[6]&r_0_addr[3],
r_2_addr[3]&r_1_addr[6]&r_0_addr[2],
r_2_addr[3]&r_1_addr[6]&r_0_addr[1],
r_2_addr[3]&r_1_addr[6]&r_0_addr[0],
r_2_addr[3]&r_1_addr[5]&r_0_addr[15],
r_2_addr[3]&r_1_addr[5]&r_0_addr[14],
r_2_addr[3]&r_1_addr[5]&r_0_addr[13],
r_2_addr[3]&r_1_addr[5]&r_0_addr[12],
r_2_addr[3]&r_1_addr[5]&r_0_addr[11],
r_2_addr[3]&r_1_addr[5]&r_0_addr[10],
r_2_addr[3]&r_1_addr[5]&r_0_addr[9],
r_2_addr[3]&r_1_addr[5]&r_0_addr[8],
r_2_addr[3]&r_1_addr[5]&r_0_addr[7],
r_2_addr[3]&r_1_addr[5]&r_0_addr[6],
r_2_addr[3]&r_1_addr[5]&r_0_addr[5],
r_2_addr[3]&r_1_addr[5]&r_0_addr[4],
r_2_addr[3]&r_1_addr[5]&r_0_addr[3],
r_2_addr[3]&r_1_addr[5]&r_0_addr[2],
r_2_addr[3]&r_1_addr[5]&r_0_addr[1],
r_2_addr[3]&r_1_addr[5]&r_0_addr[0],
r_2_addr[3]&r_1_addr[4]&r_0_addr[15],
r_2_addr[3]&r_1_addr[4]&r_0_addr[14],
r_2_addr[3]&r_1_addr[4]&r_0_addr[13],
r_2_addr[3]&r_1_addr[4]&r_0_addr[12],
r_2_addr[3]&r_1_addr[4]&r_0_addr[11],
r_2_addr[3]&r_1_addr[4]&r_0_addr[10],
r_2_addr[3]&r_1_addr[4]&r_0_addr[9],
r_2_addr[3]&r_1_addr[4]&r_0_addr[8],
r_2_addr[3]&r_1_addr[4]&r_0_addr[7],
r_2_addr[3]&r_1_addr[4]&r_0_addr[6],
r_2_addr[3]&r_1_addr[4]&r_0_addr[5],
r_2_addr[3]&r_1_addr[4]&r_0_addr[4],
r_2_addr[3]&r_1_addr[4]&r_0_addr[3],
r_2_addr[3]&r_1_addr[4]&r_0_addr[2],
r_2_addr[3]&r_1_addr[4]&r_0_addr[1],
r_2_addr[3]&r_1_addr[4]&r_0_addr[0],
r_2_addr[3]&r_1_addr[3]&r_0_addr[15],
r_2_addr[3]&r_1_addr[3]&r_0_addr[14],
r_2_addr[3]&r_1_addr[3]&r_0_addr[13],
r_2_addr[3]&r_1_addr[3]&r_0_addr[12],
r_2_addr[3]&r_1_addr[3]&r_0_addr[11],
r_2_addr[3]&r_1_addr[3]&r_0_addr[10],
r_2_addr[3]&r_1_addr[3]&r_0_addr[9],
r_2_addr[3]&r_1_addr[3]&r_0_addr[8],
r_2_addr[3]&r_1_addr[3]&r_0_addr[7],
r_2_addr[3]&r_1_addr[3]&r_0_addr[6],
r_2_addr[3]&r_1_addr[3]&r_0_addr[5],
r_2_addr[3]&r_1_addr[3]&r_0_addr[4],
r_2_addr[3]&r_1_addr[3]&r_0_addr[3],
r_2_addr[3]&r_1_addr[3]&r_0_addr[2],
r_2_addr[3]&r_1_addr[3]&r_0_addr[1],
r_2_addr[3]&r_1_addr[3]&r_0_addr[0],
r_2_addr[3]&r_1_addr[2]&r_0_addr[15],
r_2_addr[3]&r_1_addr[2]&r_0_addr[14],
r_2_addr[3]&r_1_addr[2]&r_0_addr[13],
r_2_addr[3]&r_1_addr[2]&r_0_addr[12],
r_2_addr[3]&r_1_addr[2]&r_0_addr[11],
r_2_addr[3]&r_1_addr[2]&r_0_addr[10],
r_2_addr[3]&r_1_addr[2]&r_0_addr[9],
r_2_addr[3]&r_1_addr[2]&r_0_addr[8],
r_2_addr[3]&r_1_addr[2]&r_0_addr[7],
r_2_addr[3]&r_1_addr[2]&r_0_addr[6],
r_2_addr[3]&r_1_addr[2]&r_0_addr[5],
r_2_addr[3]&r_1_addr[2]&r_0_addr[4],
r_2_addr[3]&r_1_addr[2]&r_0_addr[3],
r_2_addr[3]&r_1_addr[2]&r_0_addr[2],
r_2_addr[3]&r_1_addr[2]&r_0_addr[1],
r_2_addr[3]&r_1_addr[2]&r_0_addr[0],
r_2_addr[3]&r_1_addr[1]&r_0_addr[15],
r_2_addr[3]&r_1_addr[1]&r_0_addr[14],
r_2_addr[3]&r_1_addr[1]&r_0_addr[13],
r_2_addr[3]&r_1_addr[1]&r_0_addr[12],
r_2_addr[3]&r_1_addr[1]&r_0_addr[11],
r_2_addr[3]&r_1_addr[1]&r_0_addr[10],
r_2_addr[3]&r_1_addr[1]&r_0_addr[9],
r_2_addr[3]&r_1_addr[1]&r_0_addr[8],
r_2_addr[3]&r_1_addr[1]&r_0_addr[7],
r_2_addr[3]&r_1_addr[1]&r_0_addr[6],
r_2_addr[3]&r_1_addr[1]&r_0_addr[5],
r_2_addr[3]&r_1_addr[1]&r_0_addr[4],
r_2_addr[3]&r_1_addr[1]&r_0_addr[3],
r_2_addr[3]&r_1_addr[1]&r_0_addr[2],
r_2_addr[3]&r_1_addr[1]&r_0_addr[1],
r_2_addr[3]&r_1_addr[1]&r_0_addr[0],
r_2_addr[3]&r_1_addr[0]&r_0_addr[15],
r_2_addr[3]&r_1_addr[0]&r_0_addr[14],
r_2_addr[3]&r_1_addr[0]&r_0_addr[13],
r_2_addr[3]&r_1_addr[0]&r_0_addr[12],
r_2_addr[3]&r_1_addr[0]&r_0_addr[11],
r_2_addr[3]&r_1_addr[0]&r_0_addr[10],
r_2_addr[3]&r_1_addr[0]&r_0_addr[9],
r_2_addr[3]&r_1_addr[0]&r_0_addr[8],
r_2_addr[3]&r_1_addr[0]&r_0_addr[7],
r_2_addr[3]&r_1_addr[0]&r_0_addr[6],
r_2_addr[3]&r_1_addr[0]&r_0_addr[5],
r_2_addr[3]&r_1_addr[0]&r_0_addr[4],
r_2_addr[3]&r_1_addr[0]&r_0_addr[3],
r_2_addr[3]&r_1_addr[0]&r_0_addr[2],
r_2_addr[3]&r_1_addr[0]&r_0_addr[1],
r_2_addr[3]&r_1_addr[0]&r_0_addr[0],
r_2_addr[2]&r_1_addr[15]&r_0_addr[15],
r_2_addr[2]&r_1_addr[15]&r_0_addr[14],
r_2_addr[2]&r_1_addr[15]&r_0_addr[13],
r_2_addr[2]&r_1_addr[15]&r_0_addr[12],
r_2_addr[2]&r_1_addr[15]&r_0_addr[11],
r_2_addr[2]&r_1_addr[15]&r_0_addr[10],
r_2_addr[2]&r_1_addr[15]&r_0_addr[9],
r_2_addr[2]&r_1_addr[15]&r_0_addr[8],
r_2_addr[2]&r_1_addr[15]&r_0_addr[7],
r_2_addr[2]&r_1_addr[15]&r_0_addr[6],
r_2_addr[2]&r_1_addr[15]&r_0_addr[5],
r_2_addr[2]&r_1_addr[15]&r_0_addr[4],
r_2_addr[2]&r_1_addr[15]&r_0_addr[3],
r_2_addr[2]&r_1_addr[15]&r_0_addr[2],
r_2_addr[2]&r_1_addr[15]&r_0_addr[1],
r_2_addr[2]&r_1_addr[15]&r_0_addr[0],
r_2_addr[2]&r_1_addr[14]&r_0_addr[15],
r_2_addr[2]&r_1_addr[14]&r_0_addr[14],
r_2_addr[2]&r_1_addr[14]&r_0_addr[13],
r_2_addr[2]&r_1_addr[14]&r_0_addr[12],
r_2_addr[2]&r_1_addr[14]&r_0_addr[11],
r_2_addr[2]&r_1_addr[14]&r_0_addr[10],
r_2_addr[2]&r_1_addr[14]&r_0_addr[9],
r_2_addr[2]&r_1_addr[14]&r_0_addr[8],
r_2_addr[2]&r_1_addr[14]&r_0_addr[7],
r_2_addr[2]&r_1_addr[14]&r_0_addr[6],
r_2_addr[2]&r_1_addr[14]&r_0_addr[5],
r_2_addr[2]&r_1_addr[14]&r_0_addr[4],
r_2_addr[2]&r_1_addr[14]&r_0_addr[3],
r_2_addr[2]&r_1_addr[14]&r_0_addr[2],
r_2_addr[2]&r_1_addr[14]&r_0_addr[1],
r_2_addr[2]&r_1_addr[14]&r_0_addr[0],
r_2_addr[2]&r_1_addr[13]&r_0_addr[15],
r_2_addr[2]&r_1_addr[13]&r_0_addr[14],
r_2_addr[2]&r_1_addr[13]&r_0_addr[13],
r_2_addr[2]&r_1_addr[13]&r_0_addr[12],
r_2_addr[2]&r_1_addr[13]&r_0_addr[11],
r_2_addr[2]&r_1_addr[13]&r_0_addr[10],
r_2_addr[2]&r_1_addr[13]&r_0_addr[9],
r_2_addr[2]&r_1_addr[13]&r_0_addr[8],
r_2_addr[2]&r_1_addr[13]&r_0_addr[7],
r_2_addr[2]&r_1_addr[13]&r_0_addr[6],
r_2_addr[2]&r_1_addr[13]&r_0_addr[5],
r_2_addr[2]&r_1_addr[13]&r_0_addr[4],
r_2_addr[2]&r_1_addr[13]&r_0_addr[3],
r_2_addr[2]&r_1_addr[13]&r_0_addr[2],
r_2_addr[2]&r_1_addr[13]&r_0_addr[1],
r_2_addr[2]&r_1_addr[13]&r_0_addr[0],
r_2_addr[2]&r_1_addr[12]&r_0_addr[15],
r_2_addr[2]&r_1_addr[12]&r_0_addr[14],
r_2_addr[2]&r_1_addr[12]&r_0_addr[13],
r_2_addr[2]&r_1_addr[12]&r_0_addr[12],
r_2_addr[2]&r_1_addr[12]&r_0_addr[11],
r_2_addr[2]&r_1_addr[12]&r_0_addr[10],
r_2_addr[2]&r_1_addr[12]&r_0_addr[9],
r_2_addr[2]&r_1_addr[12]&r_0_addr[8],
r_2_addr[2]&r_1_addr[12]&r_0_addr[7],
r_2_addr[2]&r_1_addr[12]&r_0_addr[6],
r_2_addr[2]&r_1_addr[12]&r_0_addr[5],
r_2_addr[2]&r_1_addr[12]&r_0_addr[4],
r_2_addr[2]&r_1_addr[12]&r_0_addr[3],
r_2_addr[2]&r_1_addr[12]&r_0_addr[2],
r_2_addr[2]&r_1_addr[12]&r_0_addr[1],
r_2_addr[2]&r_1_addr[12]&r_0_addr[0],
r_2_addr[2]&r_1_addr[11]&r_0_addr[15],
r_2_addr[2]&r_1_addr[11]&r_0_addr[14],
r_2_addr[2]&r_1_addr[11]&r_0_addr[13],
r_2_addr[2]&r_1_addr[11]&r_0_addr[12],
r_2_addr[2]&r_1_addr[11]&r_0_addr[11],
r_2_addr[2]&r_1_addr[11]&r_0_addr[10],
r_2_addr[2]&r_1_addr[11]&r_0_addr[9],
r_2_addr[2]&r_1_addr[11]&r_0_addr[8],
r_2_addr[2]&r_1_addr[11]&r_0_addr[7],
r_2_addr[2]&r_1_addr[11]&r_0_addr[6],
r_2_addr[2]&r_1_addr[11]&r_0_addr[5],
r_2_addr[2]&r_1_addr[11]&r_0_addr[4],
r_2_addr[2]&r_1_addr[11]&r_0_addr[3],
r_2_addr[2]&r_1_addr[11]&r_0_addr[2],
r_2_addr[2]&r_1_addr[11]&r_0_addr[1],
r_2_addr[2]&r_1_addr[11]&r_0_addr[0],
r_2_addr[2]&r_1_addr[10]&r_0_addr[15],
r_2_addr[2]&r_1_addr[10]&r_0_addr[14],
r_2_addr[2]&r_1_addr[10]&r_0_addr[13],
r_2_addr[2]&r_1_addr[10]&r_0_addr[12],
r_2_addr[2]&r_1_addr[10]&r_0_addr[11],
r_2_addr[2]&r_1_addr[10]&r_0_addr[10],
r_2_addr[2]&r_1_addr[10]&r_0_addr[9],
r_2_addr[2]&r_1_addr[10]&r_0_addr[8],
r_2_addr[2]&r_1_addr[10]&r_0_addr[7],
r_2_addr[2]&r_1_addr[10]&r_0_addr[6],
r_2_addr[2]&r_1_addr[10]&r_0_addr[5],
r_2_addr[2]&r_1_addr[10]&r_0_addr[4],
r_2_addr[2]&r_1_addr[10]&r_0_addr[3],
r_2_addr[2]&r_1_addr[10]&r_0_addr[2],
r_2_addr[2]&r_1_addr[10]&r_0_addr[1],
r_2_addr[2]&r_1_addr[10]&r_0_addr[0],
r_2_addr[2]&r_1_addr[9]&r_0_addr[15],
r_2_addr[2]&r_1_addr[9]&r_0_addr[14],
r_2_addr[2]&r_1_addr[9]&r_0_addr[13],
r_2_addr[2]&r_1_addr[9]&r_0_addr[12],
r_2_addr[2]&r_1_addr[9]&r_0_addr[11],
r_2_addr[2]&r_1_addr[9]&r_0_addr[10],
r_2_addr[2]&r_1_addr[9]&r_0_addr[9],
r_2_addr[2]&r_1_addr[9]&r_0_addr[8],
r_2_addr[2]&r_1_addr[9]&r_0_addr[7],
r_2_addr[2]&r_1_addr[9]&r_0_addr[6],
r_2_addr[2]&r_1_addr[9]&r_0_addr[5],
r_2_addr[2]&r_1_addr[9]&r_0_addr[4],
r_2_addr[2]&r_1_addr[9]&r_0_addr[3],
r_2_addr[2]&r_1_addr[9]&r_0_addr[2],
r_2_addr[2]&r_1_addr[9]&r_0_addr[1],
r_2_addr[2]&r_1_addr[9]&r_0_addr[0],
r_2_addr[2]&r_1_addr[8]&r_0_addr[15],
r_2_addr[2]&r_1_addr[8]&r_0_addr[14],
r_2_addr[2]&r_1_addr[8]&r_0_addr[13],
r_2_addr[2]&r_1_addr[8]&r_0_addr[12],
r_2_addr[2]&r_1_addr[8]&r_0_addr[11],
r_2_addr[2]&r_1_addr[8]&r_0_addr[10],
r_2_addr[2]&r_1_addr[8]&r_0_addr[9],
r_2_addr[2]&r_1_addr[8]&r_0_addr[8],
r_2_addr[2]&r_1_addr[8]&r_0_addr[7],
r_2_addr[2]&r_1_addr[8]&r_0_addr[6],
r_2_addr[2]&r_1_addr[8]&r_0_addr[5],
r_2_addr[2]&r_1_addr[8]&r_0_addr[4],
r_2_addr[2]&r_1_addr[8]&r_0_addr[3],
r_2_addr[2]&r_1_addr[8]&r_0_addr[2],
r_2_addr[2]&r_1_addr[8]&r_0_addr[1],
r_2_addr[2]&r_1_addr[8]&r_0_addr[0],
r_2_addr[2]&r_1_addr[7]&r_0_addr[15],
r_2_addr[2]&r_1_addr[7]&r_0_addr[14],
r_2_addr[2]&r_1_addr[7]&r_0_addr[13],
r_2_addr[2]&r_1_addr[7]&r_0_addr[12],
r_2_addr[2]&r_1_addr[7]&r_0_addr[11],
r_2_addr[2]&r_1_addr[7]&r_0_addr[10],
r_2_addr[2]&r_1_addr[7]&r_0_addr[9],
r_2_addr[2]&r_1_addr[7]&r_0_addr[8],
r_2_addr[2]&r_1_addr[7]&r_0_addr[7],
r_2_addr[2]&r_1_addr[7]&r_0_addr[6],
r_2_addr[2]&r_1_addr[7]&r_0_addr[5],
r_2_addr[2]&r_1_addr[7]&r_0_addr[4],
r_2_addr[2]&r_1_addr[7]&r_0_addr[3],
r_2_addr[2]&r_1_addr[7]&r_0_addr[2],
r_2_addr[2]&r_1_addr[7]&r_0_addr[1],
r_2_addr[2]&r_1_addr[7]&r_0_addr[0],
r_2_addr[2]&r_1_addr[6]&r_0_addr[15],
r_2_addr[2]&r_1_addr[6]&r_0_addr[14],
r_2_addr[2]&r_1_addr[6]&r_0_addr[13],
r_2_addr[2]&r_1_addr[6]&r_0_addr[12],
r_2_addr[2]&r_1_addr[6]&r_0_addr[11],
r_2_addr[2]&r_1_addr[6]&r_0_addr[10],
r_2_addr[2]&r_1_addr[6]&r_0_addr[9],
r_2_addr[2]&r_1_addr[6]&r_0_addr[8],
r_2_addr[2]&r_1_addr[6]&r_0_addr[7],
r_2_addr[2]&r_1_addr[6]&r_0_addr[6],
r_2_addr[2]&r_1_addr[6]&r_0_addr[5],
r_2_addr[2]&r_1_addr[6]&r_0_addr[4],
r_2_addr[2]&r_1_addr[6]&r_0_addr[3],
r_2_addr[2]&r_1_addr[6]&r_0_addr[2],
r_2_addr[2]&r_1_addr[6]&r_0_addr[1],
r_2_addr[2]&r_1_addr[6]&r_0_addr[0],
r_2_addr[2]&r_1_addr[5]&r_0_addr[15],
r_2_addr[2]&r_1_addr[5]&r_0_addr[14],
r_2_addr[2]&r_1_addr[5]&r_0_addr[13],
r_2_addr[2]&r_1_addr[5]&r_0_addr[12],
r_2_addr[2]&r_1_addr[5]&r_0_addr[11],
r_2_addr[2]&r_1_addr[5]&r_0_addr[10],
r_2_addr[2]&r_1_addr[5]&r_0_addr[9],
r_2_addr[2]&r_1_addr[5]&r_0_addr[8],
r_2_addr[2]&r_1_addr[5]&r_0_addr[7],
r_2_addr[2]&r_1_addr[5]&r_0_addr[6],
r_2_addr[2]&r_1_addr[5]&r_0_addr[5],
r_2_addr[2]&r_1_addr[5]&r_0_addr[4],
r_2_addr[2]&r_1_addr[5]&r_0_addr[3],
r_2_addr[2]&r_1_addr[5]&r_0_addr[2],
r_2_addr[2]&r_1_addr[5]&r_0_addr[1],
r_2_addr[2]&r_1_addr[5]&r_0_addr[0],
r_2_addr[2]&r_1_addr[4]&r_0_addr[15],
r_2_addr[2]&r_1_addr[4]&r_0_addr[14],
r_2_addr[2]&r_1_addr[4]&r_0_addr[13],
r_2_addr[2]&r_1_addr[4]&r_0_addr[12],
r_2_addr[2]&r_1_addr[4]&r_0_addr[11],
r_2_addr[2]&r_1_addr[4]&r_0_addr[10],
r_2_addr[2]&r_1_addr[4]&r_0_addr[9],
r_2_addr[2]&r_1_addr[4]&r_0_addr[8],
r_2_addr[2]&r_1_addr[4]&r_0_addr[7],
r_2_addr[2]&r_1_addr[4]&r_0_addr[6],
r_2_addr[2]&r_1_addr[4]&r_0_addr[5],
r_2_addr[2]&r_1_addr[4]&r_0_addr[4],
r_2_addr[2]&r_1_addr[4]&r_0_addr[3],
r_2_addr[2]&r_1_addr[4]&r_0_addr[2],
r_2_addr[2]&r_1_addr[4]&r_0_addr[1],
r_2_addr[2]&r_1_addr[4]&r_0_addr[0],
r_2_addr[2]&r_1_addr[3]&r_0_addr[15],
r_2_addr[2]&r_1_addr[3]&r_0_addr[14],
r_2_addr[2]&r_1_addr[3]&r_0_addr[13],
r_2_addr[2]&r_1_addr[3]&r_0_addr[12],
r_2_addr[2]&r_1_addr[3]&r_0_addr[11],
r_2_addr[2]&r_1_addr[3]&r_0_addr[10],
r_2_addr[2]&r_1_addr[3]&r_0_addr[9],
r_2_addr[2]&r_1_addr[3]&r_0_addr[8],
r_2_addr[2]&r_1_addr[3]&r_0_addr[7],
r_2_addr[2]&r_1_addr[3]&r_0_addr[6],
r_2_addr[2]&r_1_addr[3]&r_0_addr[5],
r_2_addr[2]&r_1_addr[3]&r_0_addr[4],
r_2_addr[2]&r_1_addr[3]&r_0_addr[3],
r_2_addr[2]&r_1_addr[3]&r_0_addr[2],
r_2_addr[2]&r_1_addr[3]&r_0_addr[1],
r_2_addr[2]&r_1_addr[3]&r_0_addr[0],
r_2_addr[2]&r_1_addr[2]&r_0_addr[15],
r_2_addr[2]&r_1_addr[2]&r_0_addr[14],
r_2_addr[2]&r_1_addr[2]&r_0_addr[13],
r_2_addr[2]&r_1_addr[2]&r_0_addr[12],
r_2_addr[2]&r_1_addr[2]&r_0_addr[11],
r_2_addr[2]&r_1_addr[2]&r_0_addr[10],
r_2_addr[2]&r_1_addr[2]&r_0_addr[9],
r_2_addr[2]&r_1_addr[2]&r_0_addr[8],
r_2_addr[2]&r_1_addr[2]&r_0_addr[7],
r_2_addr[2]&r_1_addr[2]&r_0_addr[6],
r_2_addr[2]&r_1_addr[2]&r_0_addr[5],
r_2_addr[2]&r_1_addr[2]&r_0_addr[4],
r_2_addr[2]&r_1_addr[2]&r_0_addr[3],
r_2_addr[2]&r_1_addr[2]&r_0_addr[2],
r_2_addr[2]&r_1_addr[2]&r_0_addr[1],
r_2_addr[2]&r_1_addr[2]&r_0_addr[0],
r_2_addr[2]&r_1_addr[1]&r_0_addr[15],
r_2_addr[2]&r_1_addr[1]&r_0_addr[14],
r_2_addr[2]&r_1_addr[1]&r_0_addr[13],
r_2_addr[2]&r_1_addr[1]&r_0_addr[12],
r_2_addr[2]&r_1_addr[1]&r_0_addr[11],
r_2_addr[2]&r_1_addr[1]&r_0_addr[10],
r_2_addr[2]&r_1_addr[1]&r_0_addr[9],
r_2_addr[2]&r_1_addr[1]&r_0_addr[8],
r_2_addr[2]&r_1_addr[1]&r_0_addr[7],
r_2_addr[2]&r_1_addr[1]&r_0_addr[6],
r_2_addr[2]&r_1_addr[1]&r_0_addr[5],
r_2_addr[2]&r_1_addr[1]&r_0_addr[4],
r_2_addr[2]&r_1_addr[1]&r_0_addr[3],
r_2_addr[2]&r_1_addr[1]&r_0_addr[2],
r_2_addr[2]&r_1_addr[1]&r_0_addr[1],
r_2_addr[2]&r_1_addr[1]&r_0_addr[0],
r_2_addr[2]&r_1_addr[0]&r_0_addr[15],
r_2_addr[2]&r_1_addr[0]&r_0_addr[14],
r_2_addr[2]&r_1_addr[0]&r_0_addr[13],
r_2_addr[2]&r_1_addr[0]&r_0_addr[12],
r_2_addr[2]&r_1_addr[0]&r_0_addr[11],
r_2_addr[2]&r_1_addr[0]&r_0_addr[10],
r_2_addr[2]&r_1_addr[0]&r_0_addr[9],
r_2_addr[2]&r_1_addr[0]&r_0_addr[8],
r_2_addr[2]&r_1_addr[0]&r_0_addr[7],
r_2_addr[2]&r_1_addr[0]&r_0_addr[6],
r_2_addr[2]&r_1_addr[0]&r_0_addr[5],
r_2_addr[2]&r_1_addr[0]&r_0_addr[4],
r_2_addr[2]&r_1_addr[0]&r_0_addr[3],
r_2_addr[2]&r_1_addr[0]&r_0_addr[2],
r_2_addr[2]&r_1_addr[0]&r_0_addr[1],
r_2_addr[2]&r_1_addr[0]&r_0_addr[0],
r_2_addr[1]&r_1_addr[15]&r_0_addr[15],
r_2_addr[1]&r_1_addr[15]&r_0_addr[14],
r_2_addr[1]&r_1_addr[15]&r_0_addr[13],
r_2_addr[1]&r_1_addr[15]&r_0_addr[12],
r_2_addr[1]&r_1_addr[15]&r_0_addr[11],
r_2_addr[1]&r_1_addr[15]&r_0_addr[10],
r_2_addr[1]&r_1_addr[15]&r_0_addr[9],
r_2_addr[1]&r_1_addr[15]&r_0_addr[8],
r_2_addr[1]&r_1_addr[15]&r_0_addr[7],
r_2_addr[1]&r_1_addr[15]&r_0_addr[6],
r_2_addr[1]&r_1_addr[15]&r_0_addr[5],
r_2_addr[1]&r_1_addr[15]&r_0_addr[4],
r_2_addr[1]&r_1_addr[15]&r_0_addr[3],
r_2_addr[1]&r_1_addr[15]&r_0_addr[2],
r_2_addr[1]&r_1_addr[15]&r_0_addr[1],
r_2_addr[1]&r_1_addr[15]&r_0_addr[0],
r_2_addr[1]&r_1_addr[14]&r_0_addr[15],
r_2_addr[1]&r_1_addr[14]&r_0_addr[14],
r_2_addr[1]&r_1_addr[14]&r_0_addr[13],
r_2_addr[1]&r_1_addr[14]&r_0_addr[12],
r_2_addr[1]&r_1_addr[14]&r_0_addr[11],
r_2_addr[1]&r_1_addr[14]&r_0_addr[10],
r_2_addr[1]&r_1_addr[14]&r_0_addr[9],
r_2_addr[1]&r_1_addr[14]&r_0_addr[8],
r_2_addr[1]&r_1_addr[14]&r_0_addr[7],
r_2_addr[1]&r_1_addr[14]&r_0_addr[6],
r_2_addr[1]&r_1_addr[14]&r_0_addr[5],
r_2_addr[1]&r_1_addr[14]&r_0_addr[4],
r_2_addr[1]&r_1_addr[14]&r_0_addr[3],
r_2_addr[1]&r_1_addr[14]&r_0_addr[2],
r_2_addr[1]&r_1_addr[14]&r_0_addr[1],
r_2_addr[1]&r_1_addr[14]&r_0_addr[0],
r_2_addr[1]&r_1_addr[13]&r_0_addr[15],
r_2_addr[1]&r_1_addr[13]&r_0_addr[14],
r_2_addr[1]&r_1_addr[13]&r_0_addr[13],
r_2_addr[1]&r_1_addr[13]&r_0_addr[12],
r_2_addr[1]&r_1_addr[13]&r_0_addr[11],
r_2_addr[1]&r_1_addr[13]&r_0_addr[10],
r_2_addr[1]&r_1_addr[13]&r_0_addr[9],
r_2_addr[1]&r_1_addr[13]&r_0_addr[8],
r_2_addr[1]&r_1_addr[13]&r_0_addr[7],
r_2_addr[1]&r_1_addr[13]&r_0_addr[6],
r_2_addr[1]&r_1_addr[13]&r_0_addr[5],
r_2_addr[1]&r_1_addr[13]&r_0_addr[4],
r_2_addr[1]&r_1_addr[13]&r_0_addr[3],
r_2_addr[1]&r_1_addr[13]&r_0_addr[2],
r_2_addr[1]&r_1_addr[13]&r_0_addr[1],
r_2_addr[1]&r_1_addr[13]&r_0_addr[0],
r_2_addr[1]&r_1_addr[12]&r_0_addr[15],
r_2_addr[1]&r_1_addr[12]&r_0_addr[14],
r_2_addr[1]&r_1_addr[12]&r_0_addr[13],
r_2_addr[1]&r_1_addr[12]&r_0_addr[12],
r_2_addr[1]&r_1_addr[12]&r_0_addr[11],
r_2_addr[1]&r_1_addr[12]&r_0_addr[10],
r_2_addr[1]&r_1_addr[12]&r_0_addr[9],
r_2_addr[1]&r_1_addr[12]&r_0_addr[8],
r_2_addr[1]&r_1_addr[12]&r_0_addr[7],
r_2_addr[1]&r_1_addr[12]&r_0_addr[6],
r_2_addr[1]&r_1_addr[12]&r_0_addr[5],
r_2_addr[1]&r_1_addr[12]&r_0_addr[4],
r_2_addr[1]&r_1_addr[12]&r_0_addr[3],
r_2_addr[1]&r_1_addr[12]&r_0_addr[2],
r_2_addr[1]&r_1_addr[12]&r_0_addr[1],
r_2_addr[1]&r_1_addr[12]&r_0_addr[0],
r_2_addr[1]&r_1_addr[11]&r_0_addr[15],
r_2_addr[1]&r_1_addr[11]&r_0_addr[14],
r_2_addr[1]&r_1_addr[11]&r_0_addr[13],
r_2_addr[1]&r_1_addr[11]&r_0_addr[12],
r_2_addr[1]&r_1_addr[11]&r_0_addr[11],
r_2_addr[1]&r_1_addr[11]&r_0_addr[10],
r_2_addr[1]&r_1_addr[11]&r_0_addr[9],
r_2_addr[1]&r_1_addr[11]&r_0_addr[8],
r_2_addr[1]&r_1_addr[11]&r_0_addr[7],
r_2_addr[1]&r_1_addr[11]&r_0_addr[6],
r_2_addr[1]&r_1_addr[11]&r_0_addr[5],
r_2_addr[1]&r_1_addr[11]&r_0_addr[4],
r_2_addr[1]&r_1_addr[11]&r_0_addr[3],
r_2_addr[1]&r_1_addr[11]&r_0_addr[2],
r_2_addr[1]&r_1_addr[11]&r_0_addr[1],
r_2_addr[1]&r_1_addr[11]&r_0_addr[0],
r_2_addr[1]&r_1_addr[10]&r_0_addr[15],
r_2_addr[1]&r_1_addr[10]&r_0_addr[14],
r_2_addr[1]&r_1_addr[10]&r_0_addr[13],
r_2_addr[1]&r_1_addr[10]&r_0_addr[12],
r_2_addr[1]&r_1_addr[10]&r_0_addr[11],
r_2_addr[1]&r_1_addr[10]&r_0_addr[10],
r_2_addr[1]&r_1_addr[10]&r_0_addr[9],
r_2_addr[1]&r_1_addr[10]&r_0_addr[8],
r_2_addr[1]&r_1_addr[10]&r_0_addr[7],
r_2_addr[1]&r_1_addr[10]&r_0_addr[6],
r_2_addr[1]&r_1_addr[10]&r_0_addr[5],
r_2_addr[1]&r_1_addr[10]&r_0_addr[4],
r_2_addr[1]&r_1_addr[10]&r_0_addr[3],
r_2_addr[1]&r_1_addr[10]&r_0_addr[2],
r_2_addr[1]&r_1_addr[10]&r_0_addr[1],
r_2_addr[1]&r_1_addr[10]&r_0_addr[0],
r_2_addr[1]&r_1_addr[9]&r_0_addr[15],
r_2_addr[1]&r_1_addr[9]&r_0_addr[14],
r_2_addr[1]&r_1_addr[9]&r_0_addr[13],
r_2_addr[1]&r_1_addr[9]&r_0_addr[12],
r_2_addr[1]&r_1_addr[9]&r_0_addr[11],
r_2_addr[1]&r_1_addr[9]&r_0_addr[10],
r_2_addr[1]&r_1_addr[9]&r_0_addr[9],
r_2_addr[1]&r_1_addr[9]&r_0_addr[8],
r_2_addr[1]&r_1_addr[9]&r_0_addr[7],
r_2_addr[1]&r_1_addr[9]&r_0_addr[6],
r_2_addr[1]&r_1_addr[9]&r_0_addr[5],
r_2_addr[1]&r_1_addr[9]&r_0_addr[4],
r_2_addr[1]&r_1_addr[9]&r_0_addr[3],
r_2_addr[1]&r_1_addr[9]&r_0_addr[2],
r_2_addr[1]&r_1_addr[9]&r_0_addr[1],
r_2_addr[1]&r_1_addr[9]&r_0_addr[0],
r_2_addr[1]&r_1_addr[8]&r_0_addr[15],
r_2_addr[1]&r_1_addr[8]&r_0_addr[14],
r_2_addr[1]&r_1_addr[8]&r_0_addr[13],
r_2_addr[1]&r_1_addr[8]&r_0_addr[12],
r_2_addr[1]&r_1_addr[8]&r_0_addr[11],
r_2_addr[1]&r_1_addr[8]&r_0_addr[10],
r_2_addr[1]&r_1_addr[8]&r_0_addr[9],
r_2_addr[1]&r_1_addr[8]&r_0_addr[8],
r_2_addr[1]&r_1_addr[8]&r_0_addr[7],
r_2_addr[1]&r_1_addr[8]&r_0_addr[6],
r_2_addr[1]&r_1_addr[8]&r_0_addr[5],
r_2_addr[1]&r_1_addr[8]&r_0_addr[4],
r_2_addr[1]&r_1_addr[8]&r_0_addr[3],
r_2_addr[1]&r_1_addr[8]&r_0_addr[2],
r_2_addr[1]&r_1_addr[8]&r_0_addr[1],
r_2_addr[1]&r_1_addr[8]&r_0_addr[0],
r_2_addr[1]&r_1_addr[7]&r_0_addr[15],
r_2_addr[1]&r_1_addr[7]&r_0_addr[14],
r_2_addr[1]&r_1_addr[7]&r_0_addr[13],
r_2_addr[1]&r_1_addr[7]&r_0_addr[12],
r_2_addr[1]&r_1_addr[7]&r_0_addr[11],
r_2_addr[1]&r_1_addr[7]&r_0_addr[10],
r_2_addr[1]&r_1_addr[7]&r_0_addr[9],
r_2_addr[1]&r_1_addr[7]&r_0_addr[8],
r_2_addr[1]&r_1_addr[7]&r_0_addr[7],
r_2_addr[1]&r_1_addr[7]&r_0_addr[6],
r_2_addr[1]&r_1_addr[7]&r_0_addr[5],
r_2_addr[1]&r_1_addr[7]&r_0_addr[4],
r_2_addr[1]&r_1_addr[7]&r_0_addr[3],
r_2_addr[1]&r_1_addr[7]&r_0_addr[2],
r_2_addr[1]&r_1_addr[7]&r_0_addr[1],
r_2_addr[1]&r_1_addr[7]&r_0_addr[0],
r_2_addr[1]&r_1_addr[6]&r_0_addr[15],
r_2_addr[1]&r_1_addr[6]&r_0_addr[14],
r_2_addr[1]&r_1_addr[6]&r_0_addr[13],
r_2_addr[1]&r_1_addr[6]&r_0_addr[12],
r_2_addr[1]&r_1_addr[6]&r_0_addr[11],
r_2_addr[1]&r_1_addr[6]&r_0_addr[10],
r_2_addr[1]&r_1_addr[6]&r_0_addr[9],
r_2_addr[1]&r_1_addr[6]&r_0_addr[8],
r_2_addr[1]&r_1_addr[6]&r_0_addr[7],
r_2_addr[1]&r_1_addr[6]&r_0_addr[6],
r_2_addr[1]&r_1_addr[6]&r_0_addr[5],
r_2_addr[1]&r_1_addr[6]&r_0_addr[4],
r_2_addr[1]&r_1_addr[6]&r_0_addr[3],
r_2_addr[1]&r_1_addr[6]&r_0_addr[2],
r_2_addr[1]&r_1_addr[6]&r_0_addr[1],
r_2_addr[1]&r_1_addr[6]&r_0_addr[0],
r_2_addr[1]&r_1_addr[5]&r_0_addr[15],
r_2_addr[1]&r_1_addr[5]&r_0_addr[14],
r_2_addr[1]&r_1_addr[5]&r_0_addr[13],
r_2_addr[1]&r_1_addr[5]&r_0_addr[12],
r_2_addr[1]&r_1_addr[5]&r_0_addr[11],
r_2_addr[1]&r_1_addr[5]&r_0_addr[10],
r_2_addr[1]&r_1_addr[5]&r_0_addr[9],
r_2_addr[1]&r_1_addr[5]&r_0_addr[8],
r_2_addr[1]&r_1_addr[5]&r_0_addr[7],
r_2_addr[1]&r_1_addr[5]&r_0_addr[6],
r_2_addr[1]&r_1_addr[5]&r_0_addr[5],
r_2_addr[1]&r_1_addr[5]&r_0_addr[4],
r_2_addr[1]&r_1_addr[5]&r_0_addr[3],
r_2_addr[1]&r_1_addr[5]&r_0_addr[2],
r_2_addr[1]&r_1_addr[5]&r_0_addr[1],
r_2_addr[1]&r_1_addr[5]&r_0_addr[0],
r_2_addr[1]&r_1_addr[4]&r_0_addr[15],
r_2_addr[1]&r_1_addr[4]&r_0_addr[14],
r_2_addr[1]&r_1_addr[4]&r_0_addr[13],
r_2_addr[1]&r_1_addr[4]&r_0_addr[12],
r_2_addr[1]&r_1_addr[4]&r_0_addr[11],
r_2_addr[1]&r_1_addr[4]&r_0_addr[10],
r_2_addr[1]&r_1_addr[4]&r_0_addr[9],
r_2_addr[1]&r_1_addr[4]&r_0_addr[8],
r_2_addr[1]&r_1_addr[4]&r_0_addr[7],
r_2_addr[1]&r_1_addr[4]&r_0_addr[6],
r_2_addr[1]&r_1_addr[4]&r_0_addr[5],
r_2_addr[1]&r_1_addr[4]&r_0_addr[4],
r_2_addr[1]&r_1_addr[4]&r_0_addr[3],
r_2_addr[1]&r_1_addr[4]&r_0_addr[2],
r_2_addr[1]&r_1_addr[4]&r_0_addr[1],
r_2_addr[1]&r_1_addr[4]&r_0_addr[0],
r_2_addr[1]&r_1_addr[3]&r_0_addr[15],
r_2_addr[1]&r_1_addr[3]&r_0_addr[14],
r_2_addr[1]&r_1_addr[3]&r_0_addr[13],
r_2_addr[1]&r_1_addr[3]&r_0_addr[12],
r_2_addr[1]&r_1_addr[3]&r_0_addr[11],
r_2_addr[1]&r_1_addr[3]&r_0_addr[10],
r_2_addr[1]&r_1_addr[3]&r_0_addr[9],
r_2_addr[1]&r_1_addr[3]&r_0_addr[8],
r_2_addr[1]&r_1_addr[3]&r_0_addr[7],
r_2_addr[1]&r_1_addr[3]&r_0_addr[6],
r_2_addr[1]&r_1_addr[3]&r_0_addr[5],
r_2_addr[1]&r_1_addr[3]&r_0_addr[4],
r_2_addr[1]&r_1_addr[3]&r_0_addr[3],
r_2_addr[1]&r_1_addr[3]&r_0_addr[2],
r_2_addr[1]&r_1_addr[3]&r_0_addr[1],
r_2_addr[1]&r_1_addr[3]&r_0_addr[0],
r_2_addr[1]&r_1_addr[2]&r_0_addr[15],
r_2_addr[1]&r_1_addr[2]&r_0_addr[14],
r_2_addr[1]&r_1_addr[2]&r_0_addr[13],
r_2_addr[1]&r_1_addr[2]&r_0_addr[12],
r_2_addr[1]&r_1_addr[2]&r_0_addr[11],
r_2_addr[1]&r_1_addr[2]&r_0_addr[10],
r_2_addr[1]&r_1_addr[2]&r_0_addr[9],
r_2_addr[1]&r_1_addr[2]&r_0_addr[8],
r_2_addr[1]&r_1_addr[2]&r_0_addr[7],
r_2_addr[1]&r_1_addr[2]&r_0_addr[6],
r_2_addr[1]&r_1_addr[2]&r_0_addr[5],
r_2_addr[1]&r_1_addr[2]&r_0_addr[4],
r_2_addr[1]&r_1_addr[2]&r_0_addr[3],
r_2_addr[1]&r_1_addr[2]&r_0_addr[2],
r_2_addr[1]&r_1_addr[2]&r_0_addr[1],
r_2_addr[1]&r_1_addr[2]&r_0_addr[0],
r_2_addr[1]&r_1_addr[1]&r_0_addr[15],
r_2_addr[1]&r_1_addr[1]&r_0_addr[14],
r_2_addr[1]&r_1_addr[1]&r_0_addr[13],
r_2_addr[1]&r_1_addr[1]&r_0_addr[12],
r_2_addr[1]&r_1_addr[1]&r_0_addr[11],
r_2_addr[1]&r_1_addr[1]&r_0_addr[10],
r_2_addr[1]&r_1_addr[1]&r_0_addr[9],
r_2_addr[1]&r_1_addr[1]&r_0_addr[8],
r_2_addr[1]&r_1_addr[1]&r_0_addr[7],
r_2_addr[1]&r_1_addr[1]&r_0_addr[6],
r_2_addr[1]&r_1_addr[1]&r_0_addr[5],
r_2_addr[1]&r_1_addr[1]&r_0_addr[4],
r_2_addr[1]&r_1_addr[1]&r_0_addr[3],
r_2_addr[1]&r_1_addr[1]&r_0_addr[2],
r_2_addr[1]&r_1_addr[1]&r_0_addr[1],
r_2_addr[1]&r_1_addr[1]&r_0_addr[0],
r_2_addr[1]&r_1_addr[0]&r_0_addr[15],
r_2_addr[1]&r_1_addr[0]&r_0_addr[14],
r_2_addr[1]&r_1_addr[0]&r_0_addr[13],
r_2_addr[1]&r_1_addr[0]&r_0_addr[12],
r_2_addr[1]&r_1_addr[0]&r_0_addr[11],
r_2_addr[1]&r_1_addr[0]&r_0_addr[10],
r_2_addr[1]&r_1_addr[0]&r_0_addr[9],
r_2_addr[1]&r_1_addr[0]&r_0_addr[8],
r_2_addr[1]&r_1_addr[0]&r_0_addr[7],
r_2_addr[1]&r_1_addr[0]&r_0_addr[6],
r_2_addr[1]&r_1_addr[0]&r_0_addr[5],
r_2_addr[1]&r_1_addr[0]&r_0_addr[4],
r_2_addr[1]&r_1_addr[0]&r_0_addr[3],
r_2_addr[1]&r_1_addr[0]&r_0_addr[2],
r_2_addr[1]&r_1_addr[0]&r_0_addr[1],
r_2_addr[1]&r_1_addr[0]&r_0_addr[0],
r_2_addr[0]&r_1_addr[15]&r_0_addr[15],
r_2_addr[0]&r_1_addr[15]&r_0_addr[14],
r_2_addr[0]&r_1_addr[15]&r_0_addr[13],
r_2_addr[0]&r_1_addr[15]&r_0_addr[12],
r_2_addr[0]&r_1_addr[15]&r_0_addr[11],
r_2_addr[0]&r_1_addr[15]&r_0_addr[10],
r_2_addr[0]&r_1_addr[15]&r_0_addr[9],
r_2_addr[0]&r_1_addr[15]&r_0_addr[8],
r_2_addr[0]&r_1_addr[15]&r_0_addr[7],
r_2_addr[0]&r_1_addr[15]&r_0_addr[6],
r_2_addr[0]&r_1_addr[15]&r_0_addr[5],
r_2_addr[0]&r_1_addr[15]&r_0_addr[4],
r_2_addr[0]&r_1_addr[15]&r_0_addr[3],
r_2_addr[0]&r_1_addr[15]&r_0_addr[2],
r_2_addr[0]&r_1_addr[15]&r_0_addr[1],
r_2_addr[0]&r_1_addr[15]&r_0_addr[0],
r_2_addr[0]&r_1_addr[14]&r_0_addr[15],
r_2_addr[0]&r_1_addr[14]&r_0_addr[14],
r_2_addr[0]&r_1_addr[14]&r_0_addr[13],
r_2_addr[0]&r_1_addr[14]&r_0_addr[12],
r_2_addr[0]&r_1_addr[14]&r_0_addr[11],
r_2_addr[0]&r_1_addr[14]&r_0_addr[10],
r_2_addr[0]&r_1_addr[14]&r_0_addr[9],
r_2_addr[0]&r_1_addr[14]&r_0_addr[8],
r_2_addr[0]&r_1_addr[14]&r_0_addr[7],
r_2_addr[0]&r_1_addr[14]&r_0_addr[6],
r_2_addr[0]&r_1_addr[14]&r_0_addr[5],
r_2_addr[0]&r_1_addr[14]&r_0_addr[4],
r_2_addr[0]&r_1_addr[14]&r_0_addr[3],
r_2_addr[0]&r_1_addr[14]&r_0_addr[2],
r_2_addr[0]&r_1_addr[14]&r_0_addr[1],
r_2_addr[0]&r_1_addr[14]&r_0_addr[0],
r_2_addr[0]&r_1_addr[13]&r_0_addr[15],
r_2_addr[0]&r_1_addr[13]&r_0_addr[14],
r_2_addr[0]&r_1_addr[13]&r_0_addr[13],
r_2_addr[0]&r_1_addr[13]&r_0_addr[12],
r_2_addr[0]&r_1_addr[13]&r_0_addr[11],
r_2_addr[0]&r_1_addr[13]&r_0_addr[10],
r_2_addr[0]&r_1_addr[13]&r_0_addr[9],
r_2_addr[0]&r_1_addr[13]&r_0_addr[8],
r_2_addr[0]&r_1_addr[13]&r_0_addr[7],
r_2_addr[0]&r_1_addr[13]&r_0_addr[6],
r_2_addr[0]&r_1_addr[13]&r_0_addr[5],
r_2_addr[0]&r_1_addr[13]&r_0_addr[4],
r_2_addr[0]&r_1_addr[13]&r_0_addr[3],
r_2_addr[0]&r_1_addr[13]&r_0_addr[2],
r_2_addr[0]&r_1_addr[13]&r_0_addr[1],
r_2_addr[0]&r_1_addr[13]&r_0_addr[0],
r_2_addr[0]&r_1_addr[12]&r_0_addr[15],
r_2_addr[0]&r_1_addr[12]&r_0_addr[14],
r_2_addr[0]&r_1_addr[12]&r_0_addr[13],
r_2_addr[0]&r_1_addr[12]&r_0_addr[12],
r_2_addr[0]&r_1_addr[12]&r_0_addr[11],
r_2_addr[0]&r_1_addr[12]&r_0_addr[10],
r_2_addr[0]&r_1_addr[12]&r_0_addr[9],
r_2_addr[0]&r_1_addr[12]&r_0_addr[8],
r_2_addr[0]&r_1_addr[12]&r_0_addr[7],
r_2_addr[0]&r_1_addr[12]&r_0_addr[6],
r_2_addr[0]&r_1_addr[12]&r_0_addr[5],
r_2_addr[0]&r_1_addr[12]&r_0_addr[4],
r_2_addr[0]&r_1_addr[12]&r_0_addr[3],
r_2_addr[0]&r_1_addr[12]&r_0_addr[2],
r_2_addr[0]&r_1_addr[12]&r_0_addr[1],
r_2_addr[0]&r_1_addr[12]&r_0_addr[0],
r_2_addr[0]&r_1_addr[11]&r_0_addr[15],
r_2_addr[0]&r_1_addr[11]&r_0_addr[14],
r_2_addr[0]&r_1_addr[11]&r_0_addr[13],
r_2_addr[0]&r_1_addr[11]&r_0_addr[12],
r_2_addr[0]&r_1_addr[11]&r_0_addr[11],
r_2_addr[0]&r_1_addr[11]&r_0_addr[10],
r_2_addr[0]&r_1_addr[11]&r_0_addr[9],
r_2_addr[0]&r_1_addr[11]&r_0_addr[8],
r_2_addr[0]&r_1_addr[11]&r_0_addr[7],
r_2_addr[0]&r_1_addr[11]&r_0_addr[6],
r_2_addr[0]&r_1_addr[11]&r_0_addr[5],
r_2_addr[0]&r_1_addr[11]&r_0_addr[4],
r_2_addr[0]&r_1_addr[11]&r_0_addr[3],
r_2_addr[0]&r_1_addr[11]&r_0_addr[2],
r_2_addr[0]&r_1_addr[11]&r_0_addr[1],
r_2_addr[0]&r_1_addr[11]&r_0_addr[0],
r_2_addr[0]&r_1_addr[10]&r_0_addr[15],
r_2_addr[0]&r_1_addr[10]&r_0_addr[14],
r_2_addr[0]&r_1_addr[10]&r_0_addr[13],
r_2_addr[0]&r_1_addr[10]&r_0_addr[12],
r_2_addr[0]&r_1_addr[10]&r_0_addr[11],
r_2_addr[0]&r_1_addr[10]&r_0_addr[10],
r_2_addr[0]&r_1_addr[10]&r_0_addr[9],
r_2_addr[0]&r_1_addr[10]&r_0_addr[8],
r_2_addr[0]&r_1_addr[10]&r_0_addr[7],
r_2_addr[0]&r_1_addr[10]&r_0_addr[6],
r_2_addr[0]&r_1_addr[10]&r_0_addr[5],
r_2_addr[0]&r_1_addr[10]&r_0_addr[4],
r_2_addr[0]&r_1_addr[10]&r_0_addr[3],
r_2_addr[0]&r_1_addr[10]&r_0_addr[2],
r_2_addr[0]&r_1_addr[10]&r_0_addr[1],
r_2_addr[0]&r_1_addr[10]&r_0_addr[0],
r_2_addr[0]&r_1_addr[9]&r_0_addr[15],
r_2_addr[0]&r_1_addr[9]&r_0_addr[14],
r_2_addr[0]&r_1_addr[9]&r_0_addr[13],
r_2_addr[0]&r_1_addr[9]&r_0_addr[12],
r_2_addr[0]&r_1_addr[9]&r_0_addr[11],
r_2_addr[0]&r_1_addr[9]&r_0_addr[10],
r_2_addr[0]&r_1_addr[9]&r_0_addr[9],
r_2_addr[0]&r_1_addr[9]&r_0_addr[8],
r_2_addr[0]&r_1_addr[9]&r_0_addr[7],
r_2_addr[0]&r_1_addr[9]&r_0_addr[6],
r_2_addr[0]&r_1_addr[9]&r_0_addr[5],
r_2_addr[0]&r_1_addr[9]&r_0_addr[4],
r_2_addr[0]&r_1_addr[9]&r_0_addr[3],
r_2_addr[0]&r_1_addr[9]&r_0_addr[2],
r_2_addr[0]&r_1_addr[9]&r_0_addr[1],
r_2_addr[0]&r_1_addr[9]&r_0_addr[0],
r_2_addr[0]&r_1_addr[8]&r_0_addr[15],
r_2_addr[0]&r_1_addr[8]&r_0_addr[14],
r_2_addr[0]&r_1_addr[8]&r_0_addr[13],
r_2_addr[0]&r_1_addr[8]&r_0_addr[12],
r_2_addr[0]&r_1_addr[8]&r_0_addr[11],
r_2_addr[0]&r_1_addr[8]&r_0_addr[10],
r_2_addr[0]&r_1_addr[8]&r_0_addr[9],
r_2_addr[0]&r_1_addr[8]&r_0_addr[8],
r_2_addr[0]&r_1_addr[8]&r_0_addr[7],
r_2_addr[0]&r_1_addr[8]&r_0_addr[6],
r_2_addr[0]&r_1_addr[8]&r_0_addr[5],
r_2_addr[0]&r_1_addr[8]&r_0_addr[4],
r_2_addr[0]&r_1_addr[8]&r_0_addr[3],
r_2_addr[0]&r_1_addr[8]&r_0_addr[2],
r_2_addr[0]&r_1_addr[8]&r_0_addr[1],
r_2_addr[0]&r_1_addr[8]&r_0_addr[0],
r_2_addr[0]&r_1_addr[7]&r_0_addr[15],
r_2_addr[0]&r_1_addr[7]&r_0_addr[14],
r_2_addr[0]&r_1_addr[7]&r_0_addr[13],
r_2_addr[0]&r_1_addr[7]&r_0_addr[12],
r_2_addr[0]&r_1_addr[7]&r_0_addr[11],
r_2_addr[0]&r_1_addr[7]&r_0_addr[10],
r_2_addr[0]&r_1_addr[7]&r_0_addr[9],
r_2_addr[0]&r_1_addr[7]&r_0_addr[8],
r_2_addr[0]&r_1_addr[7]&r_0_addr[7],
r_2_addr[0]&r_1_addr[7]&r_0_addr[6],
r_2_addr[0]&r_1_addr[7]&r_0_addr[5],
r_2_addr[0]&r_1_addr[7]&r_0_addr[4],
r_2_addr[0]&r_1_addr[7]&r_0_addr[3],
r_2_addr[0]&r_1_addr[7]&r_0_addr[2],
r_2_addr[0]&r_1_addr[7]&r_0_addr[1],
r_2_addr[0]&r_1_addr[7]&r_0_addr[0],
r_2_addr[0]&r_1_addr[6]&r_0_addr[15],
r_2_addr[0]&r_1_addr[6]&r_0_addr[14],
r_2_addr[0]&r_1_addr[6]&r_0_addr[13],
r_2_addr[0]&r_1_addr[6]&r_0_addr[12],
r_2_addr[0]&r_1_addr[6]&r_0_addr[11],
r_2_addr[0]&r_1_addr[6]&r_0_addr[10],
r_2_addr[0]&r_1_addr[6]&r_0_addr[9],
r_2_addr[0]&r_1_addr[6]&r_0_addr[8],
r_2_addr[0]&r_1_addr[6]&r_0_addr[7],
r_2_addr[0]&r_1_addr[6]&r_0_addr[6],
r_2_addr[0]&r_1_addr[6]&r_0_addr[5],
r_2_addr[0]&r_1_addr[6]&r_0_addr[4],
r_2_addr[0]&r_1_addr[6]&r_0_addr[3],
r_2_addr[0]&r_1_addr[6]&r_0_addr[2],
r_2_addr[0]&r_1_addr[6]&r_0_addr[1],
r_2_addr[0]&r_1_addr[6]&r_0_addr[0],
r_2_addr[0]&r_1_addr[5]&r_0_addr[15],
r_2_addr[0]&r_1_addr[5]&r_0_addr[14],
r_2_addr[0]&r_1_addr[5]&r_0_addr[13],
r_2_addr[0]&r_1_addr[5]&r_0_addr[12],
r_2_addr[0]&r_1_addr[5]&r_0_addr[11],
r_2_addr[0]&r_1_addr[5]&r_0_addr[10],
r_2_addr[0]&r_1_addr[5]&r_0_addr[9],
r_2_addr[0]&r_1_addr[5]&r_0_addr[8],
r_2_addr[0]&r_1_addr[5]&r_0_addr[7],
r_2_addr[0]&r_1_addr[5]&r_0_addr[6],
r_2_addr[0]&r_1_addr[5]&r_0_addr[5],
r_2_addr[0]&r_1_addr[5]&r_0_addr[4],
r_2_addr[0]&r_1_addr[5]&r_0_addr[3],
r_2_addr[0]&r_1_addr[5]&r_0_addr[2],
r_2_addr[0]&r_1_addr[5]&r_0_addr[1],
r_2_addr[0]&r_1_addr[5]&r_0_addr[0],
r_2_addr[0]&r_1_addr[4]&r_0_addr[15],
r_2_addr[0]&r_1_addr[4]&r_0_addr[14],
r_2_addr[0]&r_1_addr[4]&r_0_addr[13],
r_2_addr[0]&r_1_addr[4]&r_0_addr[12],
r_2_addr[0]&r_1_addr[4]&r_0_addr[11],
r_2_addr[0]&r_1_addr[4]&r_0_addr[10],
r_2_addr[0]&r_1_addr[4]&r_0_addr[9],
r_2_addr[0]&r_1_addr[4]&r_0_addr[8],
r_2_addr[0]&r_1_addr[4]&r_0_addr[7],
r_2_addr[0]&r_1_addr[4]&r_0_addr[6],
r_2_addr[0]&r_1_addr[4]&r_0_addr[5],
r_2_addr[0]&r_1_addr[4]&r_0_addr[4],
r_2_addr[0]&r_1_addr[4]&r_0_addr[3],
r_2_addr[0]&r_1_addr[4]&r_0_addr[2],
r_2_addr[0]&r_1_addr[4]&r_0_addr[1],
r_2_addr[0]&r_1_addr[4]&r_0_addr[0],
r_2_addr[0]&r_1_addr[3]&r_0_addr[15],
r_2_addr[0]&r_1_addr[3]&r_0_addr[14],
r_2_addr[0]&r_1_addr[3]&r_0_addr[13],
r_2_addr[0]&r_1_addr[3]&r_0_addr[12],
r_2_addr[0]&r_1_addr[3]&r_0_addr[11],
r_2_addr[0]&r_1_addr[3]&r_0_addr[10],
r_2_addr[0]&r_1_addr[3]&r_0_addr[9],
r_2_addr[0]&r_1_addr[3]&r_0_addr[8],
r_2_addr[0]&r_1_addr[3]&r_0_addr[7],
r_2_addr[0]&r_1_addr[3]&r_0_addr[6],
r_2_addr[0]&r_1_addr[3]&r_0_addr[5],
r_2_addr[0]&r_1_addr[3]&r_0_addr[4],
r_2_addr[0]&r_1_addr[3]&r_0_addr[3],
r_2_addr[0]&r_1_addr[3]&r_0_addr[2],
r_2_addr[0]&r_1_addr[3]&r_0_addr[1],
r_2_addr[0]&r_1_addr[3]&r_0_addr[0],
r_2_addr[0]&r_1_addr[2]&r_0_addr[15],
r_2_addr[0]&r_1_addr[2]&r_0_addr[14],
r_2_addr[0]&r_1_addr[2]&r_0_addr[13],
r_2_addr[0]&r_1_addr[2]&r_0_addr[12],
r_2_addr[0]&r_1_addr[2]&r_0_addr[11],
r_2_addr[0]&r_1_addr[2]&r_0_addr[10],
r_2_addr[0]&r_1_addr[2]&r_0_addr[9],
r_2_addr[0]&r_1_addr[2]&r_0_addr[8],
r_2_addr[0]&r_1_addr[2]&r_0_addr[7],
r_2_addr[0]&r_1_addr[2]&r_0_addr[6],
r_2_addr[0]&r_1_addr[2]&r_0_addr[5],
r_2_addr[0]&r_1_addr[2]&r_0_addr[4],
r_2_addr[0]&r_1_addr[2]&r_0_addr[3],
r_2_addr[0]&r_1_addr[2]&r_0_addr[2],
r_2_addr[0]&r_1_addr[2]&r_0_addr[1],
r_2_addr[0]&r_1_addr[2]&r_0_addr[0],
r_2_addr[0]&r_1_addr[1]&r_0_addr[15],
r_2_addr[0]&r_1_addr[1]&r_0_addr[14],
r_2_addr[0]&r_1_addr[1]&r_0_addr[13],
r_2_addr[0]&r_1_addr[1]&r_0_addr[12],
r_2_addr[0]&r_1_addr[1]&r_0_addr[11],
r_2_addr[0]&r_1_addr[1]&r_0_addr[10],
r_2_addr[0]&r_1_addr[1]&r_0_addr[9],
r_2_addr[0]&r_1_addr[1]&r_0_addr[8],
r_2_addr[0]&r_1_addr[1]&r_0_addr[7],
r_2_addr[0]&r_1_addr[1]&r_0_addr[6],
r_2_addr[0]&r_1_addr[1]&r_0_addr[5],
r_2_addr[0]&r_1_addr[1]&r_0_addr[4],
r_2_addr[0]&r_1_addr[1]&r_0_addr[3],
r_2_addr[0]&r_1_addr[1]&r_0_addr[2],
r_2_addr[0]&r_1_addr[1]&r_0_addr[1],
r_2_addr[0]&r_1_addr[1]&r_0_addr[0],
r_2_addr[0]&r_1_addr[0]&r_0_addr[15],
r_2_addr[0]&r_1_addr[0]&r_0_addr[14],
r_2_addr[0]&r_1_addr[0]&r_0_addr[13],
r_2_addr[0]&r_1_addr[0]&r_0_addr[12],
r_2_addr[0]&r_1_addr[0]&r_0_addr[11],
r_2_addr[0]&r_1_addr[0]&r_0_addr[10],
r_2_addr[0]&r_1_addr[0]&r_0_addr[9],
r_2_addr[0]&r_1_addr[0]&r_0_addr[8],
r_2_addr[0]&r_1_addr[0]&r_0_addr[7],
r_2_addr[0]&r_1_addr[0]&r_0_addr[6],
r_2_addr[0]&r_1_addr[0]&r_0_addr[5],
r_2_addr[0]&r_1_addr[0]&r_0_addr[4],
r_2_addr[0]&r_1_addr[0]&r_0_addr[3],
r_2_addr[0]&r_1_addr[0]&r_0_addr[2],
r_2_addr[0]&r_1_addr[0]&r_0_addr[1],
r_2_addr[0]&r_1_addr[0]&r_0_addr[0]};


endmodule
