module Positional_encoding_16_4
(
    input wire[15:0] addr_src,
   output wire[63:0] addr_positional
);

assign addr_positional[63] = (addr_src[15:12]==4'b1111) ?1'b1:1'b0;
assign addr_positional[62] = (addr_src[15:12]==4'b1110) ?1'b1:1'b0;
assign addr_positional[61] = (addr_src[15:12]==4'b1101) ?1'b1:1'b0;
assign addr_positional[60] = (addr_src[15:12]==4'b1100) ?1'b1:1'b0;
assign addr_positional[59] = (addr_src[15:12]==4'b1011) ?1'b1:1'b0;
assign addr_positional[58] = (addr_src[15:12]==4'b1010) ?1'b1:1'b0;
assign addr_positional[57] = (addr_src[15:12]==4'b1001) ?1'b1:1'b0;
assign addr_positional[56] = (addr_src[15:12]==4'b1000) ?1'b1:1'b0;
assign addr_positional[55] = (addr_src[15:12]==4'b0111) ?1'b1:1'b0;
assign addr_positional[54] = (addr_src[15:12]==4'b0110) ?1'b1:1'b0;
assign addr_positional[53] = (addr_src[15:12]==4'b0101) ?1'b1:1'b0;
assign addr_positional[52] = (addr_src[15:12]==4'b0100) ?1'b1:1'b0;
assign addr_positional[51] = (addr_src[15:12]==4'b0011) ?1'b1:1'b0;
assign addr_positional[50] = (addr_src[15:12]==4'b0010) ?1'b1:1'b0;
assign addr_positional[49] = (addr_src[15:12]==4'b0001) ?1'b1:1'b0;
assign addr_positional[48] = (addr_src[15:12]==4'b0000) ?1'b1:1'b0;
assign addr_positional[47] = (addr_src[11:8]==4'b1111) ?1'b1:1'b0;
assign addr_positional[46] = (addr_src[11:8]==4'b1110) ?1'b1:1'b0;
assign addr_positional[45] = (addr_src[11:8]==4'b1101) ?1'b1:1'b0;
assign addr_positional[44] = (addr_src[11:8]==4'b1100) ?1'b1:1'b0;
assign addr_positional[43] = (addr_src[11:8]==4'b1011) ?1'b1:1'b0;
assign addr_positional[42] = (addr_src[11:8]==4'b1010) ?1'b1:1'b0;
assign addr_positional[41] = (addr_src[11:8]==4'b1001) ?1'b1:1'b0;
assign addr_positional[40] = (addr_src[11:8]==4'b1000) ?1'b1:1'b0;
assign addr_positional[39] = (addr_src[11:8]==4'b0111) ?1'b1:1'b0;
assign addr_positional[38] = (addr_src[11:8]==4'b0110) ?1'b1:1'b0;
assign addr_positional[37] = (addr_src[11:8]==4'b0101) ?1'b1:1'b0;
assign addr_positional[36] = (addr_src[11:8]==4'b0100) ?1'b1:1'b0;
assign addr_positional[35] = (addr_src[11:8]==4'b0011) ?1'b1:1'b0;
assign addr_positional[34] = (addr_src[11:8]==4'b0010) ?1'b1:1'b0;
assign addr_positional[33] = (addr_src[11:8]==4'b0001) ?1'b1:1'b0;
assign addr_positional[32] = (addr_src[11:8]==4'b0000) ?1'b1:1'b0;
assign addr_positional[31] = (addr_src[7:4]==4'b1111) ?1'b1:1'b0;
assign addr_positional[30] = (addr_src[7:4]==4'b1110) ?1'b1:1'b0;
assign addr_positional[29] = (addr_src[7:4]==4'b1101) ?1'b1:1'b0;
assign addr_positional[28] = (addr_src[7:4]==4'b1100) ?1'b1:1'b0;
assign addr_positional[27] = (addr_src[7:4]==4'b1011) ?1'b1:1'b0;
assign addr_positional[26] = (addr_src[7:4]==4'b1010) ?1'b1:1'b0;
assign addr_positional[25] = (addr_src[7:4]==4'b1001) ?1'b1:1'b0;
assign addr_positional[24] = (addr_src[7:4]==4'b1000) ?1'b1:1'b0;
assign addr_positional[23] = (addr_src[7:4]==4'b0111) ?1'b1:1'b0;
assign addr_positional[22] = (addr_src[7:4]==4'b0110) ?1'b1:1'b0;
assign addr_positional[21] = (addr_src[7:4]==4'b0101) ?1'b1:1'b0;
assign addr_positional[20] = (addr_src[7:4]==4'b0100) ?1'b1:1'b0;
assign addr_positional[19] = (addr_src[7:4]==4'b0011) ?1'b1:1'b0;
assign addr_positional[18] = (addr_src[7:4]==4'b0010) ?1'b1:1'b0;
assign addr_positional[17] = (addr_src[7:4]==4'b0001) ?1'b1:1'b0;
assign addr_positional[16] = (addr_src[7:4]==4'b0000) ?1'b1:1'b0;
assign addr_positional[15] = (addr_src[3:0]==4'b1111) ?1'b1:1'b0;
assign addr_positional[14] = (addr_src[3:0]==4'b1110) ?1'b1:1'b0;
assign addr_positional[13] = (addr_src[3:0]==4'b1101) ?1'b1:1'b0;
assign addr_positional[12] = (addr_src[3:0]==4'b1100) ?1'b1:1'b0;
assign addr_positional[11] = (addr_src[3:0]==4'b1011) ?1'b1:1'b0;
assign addr_positional[10] = (addr_src[3:0]==4'b1010) ?1'b1:1'b0;
assign addr_positional[9] = (addr_src[3:0]==4'b1001) ?1'b1:1'b0;
assign addr_positional[8] = (addr_src[3:0]==4'b1000) ?1'b1:1'b0;
assign addr_positional[7] = (addr_src[3:0]==4'b0111) ?1'b1:1'b0;
assign addr_positional[6] = (addr_src[3:0]==4'b0110) ?1'b1:1'b0;
assign addr_positional[5] = (addr_src[3:0]==4'b0101) ?1'b1:1'b0;
assign addr_positional[4] = (addr_src[3:0]==4'b0100) ?1'b1:1'b0;
assign addr_positional[3] = (addr_src[3:0]==4'b0011) ?1'b1:1'b0;
assign addr_positional[2] = (addr_src[3:0]==4'b0010) ?1'b1:1'b0;
assign addr_positional[1] = (addr_src[3:0]==4'b0001) ?1'b1:1'b0;
assign addr_positional[0] = (addr_src[3:0]==4'b0000) ?1'b1:1'b0;



endmodule
module address_decode_4
(
    input wire selector_enabled,
    input wire[15:0] addr_raw,
    input wire[63:0] addr_full,
   output wire[15:0] addr_selector,
    output wire[63:0] addr_remain
);

addr_remain = selector_enabled&addr_remain;
assign addr_selector[0] = selector_enabled&addr_raw[15];
assign addr_selector[1] = selector_enabled&addr_raw[14];
assign addr_selector[2] = selector_enabled&addr_raw[13];
assign addr_selector[3] = selector_enabled&addr_raw[12];
assign addr_selector[4] = selector_enabled&addr_raw[11];
assign addr_selector[5] = selector_enabled&addr_raw[10];
assign addr_selector[6] = selector_enabled&addr_raw[9];
assign addr_selector[7] = selector_enabled&addr_raw[8];
assign addr_selector[8] = selector_enabled&addr_raw[7];
assign addr_selector[9] = selector_enabled&addr_raw[6];
assign addr_selector[10] = selector_enabled&addr_raw[5];
assign addr_selector[11] = selector_enabled&addr_raw[4];
assign addr_selector[12] = selector_enabled&addr_raw[3];
assign addr_selector[13] = selector_enabled&addr_raw[2];
assign addr_selector[14] = selector_enabled&addr_raw[1];
assign addr_selector[15] = selector_enabled&addr_raw[0];


endmodule
module address_decode_16_4
(
input wire[15:0] addr_raw,
input wire selector_enabled,
output wire[65535:0] addr_selector
);

wire[63] addr_pos;
Positional_encoding_16_4 pe Positional_encoding_16_4(addr_raw, addr_pos);
wire[15:0] addr_selector0_0;
wire[15:0] addr_remain0_0;
address_decode_4 decoder_0_0 = address_decode_4(1'b1,addr_raw[63:48],addr_raw,addr_selector0_0,addr_remain0_0);


wire[15:0] addr_selector1_0;
wire[15:0] addr_remain1_0;
address_decode_4 decoder_1_0 = address_decode_4(addr_selector0_0[0],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_0,addr_remain1_0);


wire[15:0] addr_selector1_1;
wire[15:0] addr_remain1_1;
address_decode_4 decoder_1_1 = address_decode_4(addr_selector0_0[1],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_1,addr_remain1_1);


wire[15:0] addr_selector1_2;
wire[15:0] addr_remain1_2;
address_decode_4 decoder_1_2 = address_decode_4(addr_selector0_0[2],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_2,addr_remain1_2);


wire[15:0] addr_selector1_3;
wire[15:0] addr_remain1_3;
address_decode_4 decoder_1_3 = address_decode_4(addr_selector0_0[3],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_3,addr_remain1_3);


wire[15:0] addr_selector1_4;
wire[15:0] addr_remain1_4;
address_decode_4 decoder_1_4 = address_decode_4(addr_selector0_0[4],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_4,addr_remain1_4);


wire[15:0] addr_selector1_5;
wire[15:0] addr_remain1_5;
address_decode_4 decoder_1_5 = address_decode_4(addr_selector0_0[5],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_5,addr_remain1_5);


wire[15:0] addr_selector1_6;
wire[15:0] addr_remain1_6;
address_decode_4 decoder_1_6 = address_decode_4(addr_selector0_0[6],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_6,addr_remain1_6);


wire[15:0] addr_selector1_7;
wire[15:0] addr_remain1_7;
address_decode_4 decoder_1_7 = address_decode_4(addr_selector0_0[7],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_7,addr_remain1_7);


wire[15:0] addr_selector1_8;
wire[15:0] addr_remain1_8;
address_decode_4 decoder_1_8 = address_decode_4(addr_selector0_0[8],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_8,addr_remain1_8);


wire[15:0] addr_selector1_9;
wire[15:0] addr_remain1_9;
address_decode_4 decoder_1_9 = address_decode_4(addr_selector0_0[9],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_9,addr_remain1_9);


wire[15:0] addr_selector1_10;
wire[15:0] addr_remain1_10;
address_decode_4 decoder_1_10 = address_decode_4(addr_selector0_0[10],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_10,addr_remain1_10);


wire[15:0] addr_selector1_11;
wire[15:0] addr_remain1_11;
address_decode_4 decoder_1_11 = address_decode_4(addr_selector0_0[11],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_11,addr_remain1_11);


wire[15:0] addr_selector1_12;
wire[15:0] addr_remain1_12;
address_decode_4 decoder_1_12 = address_decode_4(addr_selector0_0[12],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_12,addr_remain1_12);


wire[15:0] addr_selector1_13;
wire[15:0] addr_remain1_13;
address_decode_4 decoder_1_13 = address_decode_4(addr_selector0_0[13],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_13,addr_remain1_13);


wire[15:0] addr_selector1_14;
wire[15:0] addr_remain1_14;
address_decode_4 decoder_1_14 = address_decode_4(addr_selector0_0[14],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_14,addr_remain1_14);


wire[15:0] addr_selector1_15;
wire[15:0] addr_remain1_15;
address_decode_4 decoder_1_15 = address_decode_4(addr_selector0_0[15],addr_remain0_0[47:32],addr_remain0_0,addr_selector1_15,addr_remain1_15);


wire[15:0] addr_selector2_0;
wire[15:0] addr_remain2_0;
address_decode_4 decoder_2_0 = address_decode_4(addr_selector1_0[0],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_0,addr_remain2_0);


wire[15:0] addr_selector2_1;
wire[15:0] addr_remain2_1;
address_decode_4 decoder_2_1 = address_decode_4(addr_selector1_0[1],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_1,addr_remain2_1);


wire[15:0] addr_selector2_2;
wire[15:0] addr_remain2_2;
address_decode_4 decoder_2_2 = address_decode_4(addr_selector1_0[2],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_2,addr_remain2_2);


wire[15:0] addr_selector2_3;
wire[15:0] addr_remain2_3;
address_decode_4 decoder_2_3 = address_decode_4(addr_selector1_0[3],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_3,addr_remain2_3);


wire[15:0] addr_selector2_4;
wire[15:0] addr_remain2_4;
address_decode_4 decoder_2_4 = address_decode_4(addr_selector1_0[4],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_4,addr_remain2_4);


wire[15:0] addr_selector2_5;
wire[15:0] addr_remain2_5;
address_decode_4 decoder_2_5 = address_decode_4(addr_selector1_0[5],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_5,addr_remain2_5);


wire[15:0] addr_selector2_6;
wire[15:0] addr_remain2_6;
address_decode_4 decoder_2_6 = address_decode_4(addr_selector1_0[6],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_6,addr_remain2_6);


wire[15:0] addr_selector2_7;
wire[15:0] addr_remain2_7;
address_decode_4 decoder_2_7 = address_decode_4(addr_selector1_0[7],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_7,addr_remain2_7);


wire[15:0] addr_selector2_8;
wire[15:0] addr_remain2_8;
address_decode_4 decoder_2_8 = address_decode_4(addr_selector1_0[8],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_8,addr_remain2_8);


wire[15:0] addr_selector2_9;
wire[15:0] addr_remain2_9;
address_decode_4 decoder_2_9 = address_decode_4(addr_selector1_0[9],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_9,addr_remain2_9);


wire[15:0] addr_selector2_10;
wire[15:0] addr_remain2_10;
address_decode_4 decoder_2_10 = address_decode_4(addr_selector1_0[10],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_10,addr_remain2_10);


wire[15:0] addr_selector2_11;
wire[15:0] addr_remain2_11;
address_decode_4 decoder_2_11 = address_decode_4(addr_selector1_0[11],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_11,addr_remain2_11);


wire[15:0] addr_selector2_12;
wire[15:0] addr_remain2_12;
address_decode_4 decoder_2_12 = address_decode_4(addr_selector1_0[12],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_12,addr_remain2_12);


wire[15:0] addr_selector2_13;
wire[15:0] addr_remain2_13;
address_decode_4 decoder_2_13 = address_decode_4(addr_selector1_0[13],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_13,addr_remain2_13);


wire[15:0] addr_selector2_14;
wire[15:0] addr_remain2_14;
address_decode_4 decoder_2_14 = address_decode_4(addr_selector1_0[14],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_14,addr_remain2_14);


wire[15:0] addr_selector2_15;
wire[15:0] addr_remain2_15;
address_decode_4 decoder_2_15 = address_decode_4(addr_selector1_0[15],addr_remain1_0[31:16],addr_remain1_0,addr_selector2_15,addr_remain2_15);


wire[15:0] addr_selector2_16;
wire[15:0] addr_remain2_16;
address_decode_4 decoder_2_16 = address_decode_4(addr_selector1_1[0],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_16,addr_remain2_16);


wire[15:0] addr_selector2_17;
wire[15:0] addr_remain2_17;
address_decode_4 decoder_2_17 = address_decode_4(addr_selector1_1[1],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_17,addr_remain2_17);


wire[15:0] addr_selector2_18;
wire[15:0] addr_remain2_18;
address_decode_4 decoder_2_18 = address_decode_4(addr_selector1_1[2],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_18,addr_remain2_18);


wire[15:0] addr_selector2_19;
wire[15:0] addr_remain2_19;
address_decode_4 decoder_2_19 = address_decode_4(addr_selector1_1[3],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_19,addr_remain2_19);


wire[15:0] addr_selector2_20;
wire[15:0] addr_remain2_20;
address_decode_4 decoder_2_20 = address_decode_4(addr_selector1_1[4],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_20,addr_remain2_20);


wire[15:0] addr_selector2_21;
wire[15:0] addr_remain2_21;
address_decode_4 decoder_2_21 = address_decode_4(addr_selector1_1[5],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_21,addr_remain2_21);


wire[15:0] addr_selector2_22;
wire[15:0] addr_remain2_22;
address_decode_4 decoder_2_22 = address_decode_4(addr_selector1_1[6],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_22,addr_remain2_22);


wire[15:0] addr_selector2_23;
wire[15:0] addr_remain2_23;
address_decode_4 decoder_2_23 = address_decode_4(addr_selector1_1[7],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_23,addr_remain2_23);


wire[15:0] addr_selector2_24;
wire[15:0] addr_remain2_24;
address_decode_4 decoder_2_24 = address_decode_4(addr_selector1_1[8],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_24,addr_remain2_24);


wire[15:0] addr_selector2_25;
wire[15:0] addr_remain2_25;
address_decode_4 decoder_2_25 = address_decode_4(addr_selector1_1[9],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_25,addr_remain2_25);


wire[15:0] addr_selector2_26;
wire[15:0] addr_remain2_26;
address_decode_4 decoder_2_26 = address_decode_4(addr_selector1_1[10],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_26,addr_remain2_26);


wire[15:0] addr_selector2_27;
wire[15:0] addr_remain2_27;
address_decode_4 decoder_2_27 = address_decode_4(addr_selector1_1[11],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_27,addr_remain2_27);


wire[15:0] addr_selector2_28;
wire[15:0] addr_remain2_28;
address_decode_4 decoder_2_28 = address_decode_4(addr_selector1_1[12],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_28,addr_remain2_28);


wire[15:0] addr_selector2_29;
wire[15:0] addr_remain2_29;
address_decode_4 decoder_2_29 = address_decode_4(addr_selector1_1[13],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_29,addr_remain2_29);


wire[15:0] addr_selector2_30;
wire[15:0] addr_remain2_30;
address_decode_4 decoder_2_30 = address_decode_4(addr_selector1_1[14],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_30,addr_remain2_30);


wire[15:0] addr_selector2_31;
wire[15:0] addr_remain2_31;
address_decode_4 decoder_2_31 = address_decode_4(addr_selector1_1[15],addr_remain1_1[31:16],addr_remain1_1,addr_selector2_31,addr_remain2_31);


wire[15:0] addr_selector2_32;
wire[15:0] addr_remain2_32;
address_decode_4 decoder_2_32 = address_decode_4(addr_selector1_2[0],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_32,addr_remain2_32);


wire[15:0] addr_selector2_33;
wire[15:0] addr_remain2_33;
address_decode_4 decoder_2_33 = address_decode_4(addr_selector1_2[1],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_33,addr_remain2_33);


wire[15:0] addr_selector2_34;
wire[15:0] addr_remain2_34;
address_decode_4 decoder_2_34 = address_decode_4(addr_selector1_2[2],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_34,addr_remain2_34);


wire[15:0] addr_selector2_35;
wire[15:0] addr_remain2_35;
address_decode_4 decoder_2_35 = address_decode_4(addr_selector1_2[3],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_35,addr_remain2_35);


wire[15:0] addr_selector2_36;
wire[15:0] addr_remain2_36;
address_decode_4 decoder_2_36 = address_decode_4(addr_selector1_2[4],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_36,addr_remain2_36);


wire[15:0] addr_selector2_37;
wire[15:0] addr_remain2_37;
address_decode_4 decoder_2_37 = address_decode_4(addr_selector1_2[5],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_37,addr_remain2_37);


wire[15:0] addr_selector2_38;
wire[15:0] addr_remain2_38;
address_decode_4 decoder_2_38 = address_decode_4(addr_selector1_2[6],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_38,addr_remain2_38);


wire[15:0] addr_selector2_39;
wire[15:0] addr_remain2_39;
address_decode_4 decoder_2_39 = address_decode_4(addr_selector1_2[7],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_39,addr_remain2_39);


wire[15:0] addr_selector2_40;
wire[15:0] addr_remain2_40;
address_decode_4 decoder_2_40 = address_decode_4(addr_selector1_2[8],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_40,addr_remain2_40);


wire[15:0] addr_selector2_41;
wire[15:0] addr_remain2_41;
address_decode_4 decoder_2_41 = address_decode_4(addr_selector1_2[9],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_41,addr_remain2_41);


wire[15:0] addr_selector2_42;
wire[15:0] addr_remain2_42;
address_decode_4 decoder_2_42 = address_decode_4(addr_selector1_2[10],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_42,addr_remain2_42);


wire[15:0] addr_selector2_43;
wire[15:0] addr_remain2_43;
address_decode_4 decoder_2_43 = address_decode_4(addr_selector1_2[11],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_43,addr_remain2_43);


wire[15:0] addr_selector2_44;
wire[15:0] addr_remain2_44;
address_decode_4 decoder_2_44 = address_decode_4(addr_selector1_2[12],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_44,addr_remain2_44);


wire[15:0] addr_selector2_45;
wire[15:0] addr_remain2_45;
address_decode_4 decoder_2_45 = address_decode_4(addr_selector1_2[13],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_45,addr_remain2_45);


wire[15:0] addr_selector2_46;
wire[15:0] addr_remain2_46;
address_decode_4 decoder_2_46 = address_decode_4(addr_selector1_2[14],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_46,addr_remain2_46);


wire[15:0] addr_selector2_47;
wire[15:0] addr_remain2_47;
address_decode_4 decoder_2_47 = address_decode_4(addr_selector1_2[15],addr_remain1_2[31:16],addr_remain1_2,addr_selector2_47,addr_remain2_47);


wire[15:0] addr_selector2_48;
wire[15:0] addr_remain2_48;
address_decode_4 decoder_2_48 = address_decode_4(addr_selector1_3[0],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_48,addr_remain2_48);


wire[15:0] addr_selector2_49;
wire[15:0] addr_remain2_49;
address_decode_4 decoder_2_49 = address_decode_4(addr_selector1_3[1],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_49,addr_remain2_49);


wire[15:0] addr_selector2_50;
wire[15:0] addr_remain2_50;
address_decode_4 decoder_2_50 = address_decode_4(addr_selector1_3[2],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_50,addr_remain2_50);


wire[15:0] addr_selector2_51;
wire[15:0] addr_remain2_51;
address_decode_4 decoder_2_51 = address_decode_4(addr_selector1_3[3],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_51,addr_remain2_51);


wire[15:0] addr_selector2_52;
wire[15:0] addr_remain2_52;
address_decode_4 decoder_2_52 = address_decode_4(addr_selector1_3[4],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_52,addr_remain2_52);


wire[15:0] addr_selector2_53;
wire[15:0] addr_remain2_53;
address_decode_4 decoder_2_53 = address_decode_4(addr_selector1_3[5],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_53,addr_remain2_53);


wire[15:0] addr_selector2_54;
wire[15:0] addr_remain2_54;
address_decode_4 decoder_2_54 = address_decode_4(addr_selector1_3[6],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_54,addr_remain2_54);


wire[15:0] addr_selector2_55;
wire[15:0] addr_remain2_55;
address_decode_4 decoder_2_55 = address_decode_4(addr_selector1_3[7],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_55,addr_remain2_55);


wire[15:0] addr_selector2_56;
wire[15:0] addr_remain2_56;
address_decode_4 decoder_2_56 = address_decode_4(addr_selector1_3[8],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_56,addr_remain2_56);


wire[15:0] addr_selector2_57;
wire[15:0] addr_remain2_57;
address_decode_4 decoder_2_57 = address_decode_4(addr_selector1_3[9],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_57,addr_remain2_57);


wire[15:0] addr_selector2_58;
wire[15:0] addr_remain2_58;
address_decode_4 decoder_2_58 = address_decode_4(addr_selector1_3[10],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_58,addr_remain2_58);


wire[15:0] addr_selector2_59;
wire[15:0] addr_remain2_59;
address_decode_4 decoder_2_59 = address_decode_4(addr_selector1_3[11],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_59,addr_remain2_59);


wire[15:0] addr_selector2_60;
wire[15:0] addr_remain2_60;
address_decode_4 decoder_2_60 = address_decode_4(addr_selector1_3[12],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_60,addr_remain2_60);


wire[15:0] addr_selector2_61;
wire[15:0] addr_remain2_61;
address_decode_4 decoder_2_61 = address_decode_4(addr_selector1_3[13],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_61,addr_remain2_61);


wire[15:0] addr_selector2_62;
wire[15:0] addr_remain2_62;
address_decode_4 decoder_2_62 = address_decode_4(addr_selector1_3[14],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_62,addr_remain2_62);


wire[15:0] addr_selector2_63;
wire[15:0] addr_remain2_63;
address_decode_4 decoder_2_63 = address_decode_4(addr_selector1_3[15],addr_remain1_3[31:16],addr_remain1_3,addr_selector2_63,addr_remain2_63);


wire[15:0] addr_selector2_64;
wire[15:0] addr_remain2_64;
address_decode_4 decoder_2_64 = address_decode_4(addr_selector1_4[0],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_64,addr_remain2_64);


wire[15:0] addr_selector2_65;
wire[15:0] addr_remain2_65;
address_decode_4 decoder_2_65 = address_decode_4(addr_selector1_4[1],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_65,addr_remain2_65);


wire[15:0] addr_selector2_66;
wire[15:0] addr_remain2_66;
address_decode_4 decoder_2_66 = address_decode_4(addr_selector1_4[2],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_66,addr_remain2_66);


wire[15:0] addr_selector2_67;
wire[15:0] addr_remain2_67;
address_decode_4 decoder_2_67 = address_decode_4(addr_selector1_4[3],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_67,addr_remain2_67);


wire[15:0] addr_selector2_68;
wire[15:0] addr_remain2_68;
address_decode_4 decoder_2_68 = address_decode_4(addr_selector1_4[4],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_68,addr_remain2_68);


wire[15:0] addr_selector2_69;
wire[15:0] addr_remain2_69;
address_decode_4 decoder_2_69 = address_decode_4(addr_selector1_4[5],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_69,addr_remain2_69);


wire[15:0] addr_selector2_70;
wire[15:0] addr_remain2_70;
address_decode_4 decoder_2_70 = address_decode_4(addr_selector1_4[6],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_70,addr_remain2_70);


wire[15:0] addr_selector2_71;
wire[15:0] addr_remain2_71;
address_decode_4 decoder_2_71 = address_decode_4(addr_selector1_4[7],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_71,addr_remain2_71);


wire[15:0] addr_selector2_72;
wire[15:0] addr_remain2_72;
address_decode_4 decoder_2_72 = address_decode_4(addr_selector1_4[8],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_72,addr_remain2_72);


wire[15:0] addr_selector2_73;
wire[15:0] addr_remain2_73;
address_decode_4 decoder_2_73 = address_decode_4(addr_selector1_4[9],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_73,addr_remain2_73);


wire[15:0] addr_selector2_74;
wire[15:0] addr_remain2_74;
address_decode_4 decoder_2_74 = address_decode_4(addr_selector1_4[10],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_74,addr_remain2_74);


wire[15:0] addr_selector2_75;
wire[15:0] addr_remain2_75;
address_decode_4 decoder_2_75 = address_decode_4(addr_selector1_4[11],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_75,addr_remain2_75);


wire[15:0] addr_selector2_76;
wire[15:0] addr_remain2_76;
address_decode_4 decoder_2_76 = address_decode_4(addr_selector1_4[12],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_76,addr_remain2_76);


wire[15:0] addr_selector2_77;
wire[15:0] addr_remain2_77;
address_decode_4 decoder_2_77 = address_decode_4(addr_selector1_4[13],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_77,addr_remain2_77);


wire[15:0] addr_selector2_78;
wire[15:0] addr_remain2_78;
address_decode_4 decoder_2_78 = address_decode_4(addr_selector1_4[14],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_78,addr_remain2_78);


wire[15:0] addr_selector2_79;
wire[15:0] addr_remain2_79;
address_decode_4 decoder_2_79 = address_decode_4(addr_selector1_4[15],addr_remain1_4[31:16],addr_remain1_4,addr_selector2_79,addr_remain2_79);


wire[15:0] addr_selector2_80;
wire[15:0] addr_remain2_80;
address_decode_4 decoder_2_80 = address_decode_4(addr_selector1_5[0],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_80,addr_remain2_80);


wire[15:0] addr_selector2_81;
wire[15:0] addr_remain2_81;
address_decode_4 decoder_2_81 = address_decode_4(addr_selector1_5[1],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_81,addr_remain2_81);


wire[15:0] addr_selector2_82;
wire[15:0] addr_remain2_82;
address_decode_4 decoder_2_82 = address_decode_4(addr_selector1_5[2],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_82,addr_remain2_82);


wire[15:0] addr_selector2_83;
wire[15:0] addr_remain2_83;
address_decode_4 decoder_2_83 = address_decode_4(addr_selector1_5[3],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_83,addr_remain2_83);


wire[15:0] addr_selector2_84;
wire[15:0] addr_remain2_84;
address_decode_4 decoder_2_84 = address_decode_4(addr_selector1_5[4],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_84,addr_remain2_84);


wire[15:0] addr_selector2_85;
wire[15:0] addr_remain2_85;
address_decode_4 decoder_2_85 = address_decode_4(addr_selector1_5[5],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_85,addr_remain2_85);


wire[15:0] addr_selector2_86;
wire[15:0] addr_remain2_86;
address_decode_4 decoder_2_86 = address_decode_4(addr_selector1_5[6],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_86,addr_remain2_86);


wire[15:0] addr_selector2_87;
wire[15:0] addr_remain2_87;
address_decode_4 decoder_2_87 = address_decode_4(addr_selector1_5[7],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_87,addr_remain2_87);


wire[15:0] addr_selector2_88;
wire[15:0] addr_remain2_88;
address_decode_4 decoder_2_88 = address_decode_4(addr_selector1_5[8],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_88,addr_remain2_88);


wire[15:0] addr_selector2_89;
wire[15:0] addr_remain2_89;
address_decode_4 decoder_2_89 = address_decode_4(addr_selector1_5[9],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_89,addr_remain2_89);


wire[15:0] addr_selector2_90;
wire[15:0] addr_remain2_90;
address_decode_4 decoder_2_90 = address_decode_4(addr_selector1_5[10],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_90,addr_remain2_90);


wire[15:0] addr_selector2_91;
wire[15:0] addr_remain2_91;
address_decode_4 decoder_2_91 = address_decode_4(addr_selector1_5[11],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_91,addr_remain2_91);


wire[15:0] addr_selector2_92;
wire[15:0] addr_remain2_92;
address_decode_4 decoder_2_92 = address_decode_4(addr_selector1_5[12],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_92,addr_remain2_92);


wire[15:0] addr_selector2_93;
wire[15:0] addr_remain2_93;
address_decode_4 decoder_2_93 = address_decode_4(addr_selector1_5[13],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_93,addr_remain2_93);


wire[15:0] addr_selector2_94;
wire[15:0] addr_remain2_94;
address_decode_4 decoder_2_94 = address_decode_4(addr_selector1_5[14],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_94,addr_remain2_94);


wire[15:0] addr_selector2_95;
wire[15:0] addr_remain2_95;
address_decode_4 decoder_2_95 = address_decode_4(addr_selector1_5[15],addr_remain1_5[31:16],addr_remain1_5,addr_selector2_95,addr_remain2_95);


wire[15:0] addr_selector2_96;
wire[15:0] addr_remain2_96;
address_decode_4 decoder_2_96 = address_decode_4(addr_selector1_6[0],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_96,addr_remain2_96);


wire[15:0] addr_selector2_97;
wire[15:0] addr_remain2_97;
address_decode_4 decoder_2_97 = address_decode_4(addr_selector1_6[1],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_97,addr_remain2_97);


wire[15:0] addr_selector2_98;
wire[15:0] addr_remain2_98;
address_decode_4 decoder_2_98 = address_decode_4(addr_selector1_6[2],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_98,addr_remain2_98);


wire[15:0] addr_selector2_99;
wire[15:0] addr_remain2_99;
address_decode_4 decoder_2_99 = address_decode_4(addr_selector1_6[3],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_99,addr_remain2_99);


wire[15:0] addr_selector2_100;
wire[15:0] addr_remain2_100;
address_decode_4 decoder_2_100 = address_decode_4(addr_selector1_6[4],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_100,addr_remain2_100);


wire[15:0] addr_selector2_101;
wire[15:0] addr_remain2_101;
address_decode_4 decoder_2_101 = address_decode_4(addr_selector1_6[5],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_101,addr_remain2_101);


wire[15:0] addr_selector2_102;
wire[15:0] addr_remain2_102;
address_decode_4 decoder_2_102 = address_decode_4(addr_selector1_6[6],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_102,addr_remain2_102);


wire[15:0] addr_selector2_103;
wire[15:0] addr_remain2_103;
address_decode_4 decoder_2_103 = address_decode_4(addr_selector1_6[7],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_103,addr_remain2_103);


wire[15:0] addr_selector2_104;
wire[15:0] addr_remain2_104;
address_decode_4 decoder_2_104 = address_decode_4(addr_selector1_6[8],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_104,addr_remain2_104);


wire[15:0] addr_selector2_105;
wire[15:0] addr_remain2_105;
address_decode_4 decoder_2_105 = address_decode_4(addr_selector1_6[9],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_105,addr_remain2_105);


wire[15:0] addr_selector2_106;
wire[15:0] addr_remain2_106;
address_decode_4 decoder_2_106 = address_decode_4(addr_selector1_6[10],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_106,addr_remain2_106);


wire[15:0] addr_selector2_107;
wire[15:0] addr_remain2_107;
address_decode_4 decoder_2_107 = address_decode_4(addr_selector1_6[11],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_107,addr_remain2_107);


wire[15:0] addr_selector2_108;
wire[15:0] addr_remain2_108;
address_decode_4 decoder_2_108 = address_decode_4(addr_selector1_6[12],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_108,addr_remain2_108);


wire[15:0] addr_selector2_109;
wire[15:0] addr_remain2_109;
address_decode_4 decoder_2_109 = address_decode_4(addr_selector1_6[13],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_109,addr_remain2_109);


wire[15:0] addr_selector2_110;
wire[15:0] addr_remain2_110;
address_decode_4 decoder_2_110 = address_decode_4(addr_selector1_6[14],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_110,addr_remain2_110);


wire[15:0] addr_selector2_111;
wire[15:0] addr_remain2_111;
address_decode_4 decoder_2_111 = address_decode_4(addr_selector1_6[15],addr_remain1_6[31:16],addr_remain1_6,addr_selector2_111,addr_remain2_111);


wire[15:0] addr_selector2_112;
wire[15:0] addr_remain2_112;
address_decode_4 decoder_2_112 = address_decode_4(addr_selector1_7[0],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_112,addr_remain2_112);


wire[15:0] addr_selector2_113;
wire[15:0] addr_remain2_113;
address_decode_4 decoder_2_113 = address_decode_4(addr_selector1_7[1],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_113,addr_remain2_113);


wire[15:0] addr_selector2_114;
wire[15:0] addr_remain2_114;
address_decode_4 decoder_2_114 = address_decode_4(addr_selector1_7[2],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_114,addr_remain2_114);


wire[15:0] addr_selector2_115;
wire[15:0] addr_remain2_115;
address_decode_4 decoder_2_115 = address_decode_4(addr_selector1_7[3],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_115,addr_remain2_115);


wire[15:0] addr_selector2_116;
wire[15:0] addr_remain2_116;
address_decode_4 decoder_2_116 = address_decode_4(addr_selector1_7[4],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_116,addr_remain2_116);


wire[15:0] addr_selector2_117;
wire[15:0] addr_remain2_117;
address_decode_4 decoder_2_117 = address_decode_4(addr_selector1_7[5],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_117,addr_remain2_117);


wire[15:0] addr_selector2_118;
wire[15:0] addr_remain2_118;
address_decode_4 decoder_2_118 = address_decode_4(addr_selector1_7[6],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_118,addr_remain2_118);


wire[15:0] addr_selector2_119;
wire[15:0] addr_remain2_119;
address_decode_4 decoder_2_119 = address_decode_4(addr_selector1_7[7],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_119,addr_remain2_119);


wire[15:0] addr_selector2_120;
wire[15:0] addr_remain2_120;
address_decode_4 decoder_2_120 = address_decode_4(addr_selector1_7[8],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_120,addr_remain2_120);


wire[15:0] addr_selector2_121;
wire[15:0] addr_remain2_121;
address_decode_4 decoder_2_121 = address_decode_4(addr_selector1_7[9],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_121,addr_remain2_121);


wire[15:0] addr_selector2_122;
wire[15:0] addr_remain2_122;
address_decode_4 decoder_2_122 = address_decode_4(addr_selector1_7[10],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_122,addr_remain2_122);


wire[15:0] addr_selector2_123;
wire[15:0] addr_remain2_123;
address_decode_4 decoder_2_123 = address_decode_4(addr_selector1_7[11],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_123,addr_remain2_123);


wire[15:0] addr_selector2_124;
wire[15:0] addr_remain2_124;
address_decode_4 decoder_2_124 = address_decode_4(addr_selector1_7[12],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_124,addr_remain2_124);


wire[15:0] addr_selector2_125;
wire[15:0] addr_remain2_125;
address_decode_4 decoder_2_125 = address_decode_4(addr_selector1_7[13],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_125,addr_remain2_125);


wire[15:0] addr_selector2_126;
wire[15:0] addr_remain2_126;
address_decode_4 decoder_2_126 = address_decode_4(addr_selector1_7[14],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_126,addr_remain2_126);


wire[15:0] addr_selector2_127;
wire[15:0] addr_remain2_127;
address_decode_4 decoder_2_127 = address_decode_4(addr_selector1_7[15],addr_remain1_7[31:16],addr_remain1_7,addr_selector2_127,addr_remain2_127);


wire[15:0] addr_selector2_128;
wire[15:0] addr_remain2_128;
address_decode_4 decoder_2_128 = address_decode_4(addr_selector1_8[0],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_128,addr_remain2_128);


wire[15:0] addr_selector2_129;
wire[15:0] addr_remain2_129;
address_decode_4 decoder_2_129 = address_decode_4(addr_selector1_8[1],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_129,addr_remain2_129);


wire[15:0] addr_selector2_130;
wire[15:0] addr_remain2_130;
address_decode_4 decoder_2_130 = address_decode_4(addr_selector1_8[2],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_130,addr_remain2_130);


wire[15:0] addr_selector2_131;
wire[15:0] addr_remain2_131;
address_decode_4 decoder_2_131 = address_decode_4(addr_selector1_8[3],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_131,addr_remain2_131);


wire[15:0] addr_selector2_132;
wire[15:0] addr_remain2_132;
address_decode_4 decoder_2_132 = address_decode_4(addr_selector1_8[4],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_132,addr_remain2_132);


wire[15:0] addr_selector2_133;
wire[15:0] addr_remain2_133;
address_decode_4 decoder_2_133 = address_decode_4(addr_selector1_8[5],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_133,addr_remain2_133);


wire[15:0] addr_selector2_134;
wire[15:0] addr_remain2_134;
address_decode_4 decoder_2_134 = address_decode_4(addr_selector1_8[6],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_134,addr_remain2_134);


wire[15:0] addr_selector2_135;
wire[15:0] addr_remain2_135;
address_decode_4 decoder_2_135 = address_decode_4(addr_selector1_8[7],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_135,addr_remain2_135);


wire[15:0] addr_selector2_136;
wire[15:0] addr_remain2_136;
address_decode_4 decoder_2_136 = address_decode_4(addr_selector1_8[8],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_136,addr_remain2_136);


wire[15:0] addr_selector2_137;
wire[15:0] addr_remain2_137;
address_decode_4 decoder_2_137 = address_decode_4(addr_selector1_8[9],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_137,addr_remain2_137);


wire[15:0] addr_selector2_138;
wire[15:0] addr_remain2_138;
address_decode_4 decoder_2_138 = address_decode_4(addr_selector1_8[10],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_138,addr_remain2_138);


wire[15:0] addr_selector2_139;
wire[15:0] addr_remain2_139;
address_decode_4 decoder_2_139 = address_decode_4(addr_selector1_8[11],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_139,addr_remain2_139);


wire[15:0] addr_selector2_140;
wire[15:0] addr_remain2_140;
address_decode_4 decoder_2_140 = address_decode_4(addr_selector1_8[12],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_140,addr_remain2_140);


wire[15:0] addr_selector2_141;
wire[15:0] addr_remain2_141;
address_decode_4 decoder_2_141 = address_decode_4(addr_selector1_8[13],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_141,addr_remain2_141);


wire[15:0] addr_selector2_142;
wire[15:0] addr_remain2_142;
address_decode_4 decoder_2_142 = address_decode_4(addr_selector1_8[14],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_142,addr_remain2_142);


wire[15:0] addr_selector2_143;
wire[15:0] addr_remain2_143;
address_decode_4 decoder_2_143 = address_decode_4(addr_selector1_8[15],addr_remain1_8[31:16],addr_remain1_8,addr_selector2_143,addr_remain2_143);


wire[15:0] addr_selector2_144;
wire[15:0] addr_remain2_144;
address_decode_4 decoder_2_144 = address_decode_4(addr_selector1_9[0],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_144,addr_remain2_144);


wire[15:0] addr_selector2_145;
wire[15:0] addr_remain2_145;
address_decode_4 decoder_2_145 = address_decode_4(addr_selector1_9[1],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_145,addr_remain2_145);


wire[15:0] addr_selector2_146;
wire[15:0] addr_remain2_146;
address_decode_4 decoder_2_146 = address_decode_4(addr_selector1_9[2],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_146,addr_remain2_146);


wire[15:0] addr_selector2_147;
wire[15:0] addr_remain2_147;
address_decode_4 decoder_2_147 = address_decode_4(addr_selector1_9[3],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_147,addr_remain2_147);


wire[15:0] addr_selector2_148;
wire[15:0] addr_remain2_148;
address_decode_4 decoder_2_148 = address_decode_4(addr_selector1_9[4],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_148,addr_remain2_148);


wire[15:0] addr_selector2_149;
wire[15:0] addr_remain2_149;
address_decode_4 decoder_2_149 = address_decode_4(addr_selector1_9[5],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_149,addr_remain2_149);


wire[15:0] addr_selector2_150;
wire[15:0] addr_remain2_150;
address_decode_4 decoder_2_150 = address_decode_4(addr_selector1_9[6],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_150,addr_remain2_150);


wire[15:0] addr_selector2_151;
wire[15:0] addr_remain2_151;
address_decode_4 decoder_2_151 = address_decode_4(addr_selector1_9[7],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_151,addr_remain2_151);


wire[15:0] addr_selector2_152;
wire[15:0] addr_remain2_152;
address_decode_4 decoder_2_152 = address_decode_4(addr_selector1_9[8],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_152,addr_remain2_152);


wire[15:0] addr_selector2_153;
wire[15:0] addr_remain2_153;
address_decode_4 decoder_2_153 = address_decode_4(addr_selector1_9[9],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_153,addr_remain2_153);


wire[15:0] addr_selector2_154;
wire[15:0] addr_remain2_154;
address_decode_4 decoder_2_154 = address_decode_4(addr_selector1_9[10],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_154,addr_remain2_154);


wire[15:0] addr_selector2_155;
wire[15:0] addr_remain2_155;
address_decode_4 decoder_2_155 = address_decode_4(addr_selector1_9[11],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_155,addr_remain2_155);


wire[15:0] addr_selector2_156;
wire[15:0] addr_remain2_156;
address_decode_4 decoder_2_156 = address_decode_4(addr_selector1_9[12],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_156,addr_remain2_156);


wire[15:0] addr_selector2_157;
wire[15:0] addr_remain2_157;
address_decode_4 decoder_2_157 = address_decode_4(addr_selector1_9[13],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_157,addr_remain2_157);


wire[15:0] addr_selector2_158;
wire[15:0] addr_remain2_158;
address_decode_4 decoder_2_158 = address_decode_4(addr_selector1_9[14],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_158,addr_remain2_158);


wire[15:0] addr_selector2_159;
wire[15:0] addr_remain2_159;
address_decode_4 decoder_2_159 = address_decode_4(addr_selector1_9[15],addr_remain1_9[31:16],addr_remain1_9,addr_selector2_159,addr_remain2_159);


wire[15:0] addr_selector2_160;
wire[15:0] addr_remain2_160;
address_decode_4 decoder_2_160 = address_decode_4(addr_selector1_10[0],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_160,addr_remain2_160);


wire[15:0] addr_selector2_161;
wire[15:0] addr_remain2_161;
address_decode_4 decoder_2_161 = address_decode_4(addr_selector1_10[1],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_161,addr_remain2_161);


wire[15:0] addr_selector2_162;
wire[15:0] addr_remain2_162;
address_decode_4 decoder_2_162 = address_decode_4(addr_selector1_10[2],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_162,addr_remain2_162);


wire[15:0] addr_selector2_163;
wire[15:0] addr_remain2_163;
address_decode_4 decoder_2_163 = address_decode_4(addr_selector1_10[3],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_163,addr_remain2_163);


wire[15:0] addr_selector2_164;
wire[15:0] addr_remain2_164;
address_decode_4 decoder_2_164 = address_decode_4(addr_selector1_10[4],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_164,addr_remain2_164);


wire[15:0] addr_selector2_165;
wire[15:0] addr_remain2_165;
address_decode_4 decoder_2_165 = address_decode_4(addr_selector1_10[5],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_165,addr_remain2_165);


wire[15:0] addr_selector2_166;
wire[15:0] addr_remain2_166;
address_decode_4 decoder_2_166 = address_decode_4(addr_selector1_10[6],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_166,addr_remain2_166);


wire[15:0] addr_selector2_167;
wire[15:0] addr_remain2_167;
address_decode_4 decoder_2_167 = address_decode_4(addr_selector1_10[7],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_167,addr_remain2_167);


wire[15:0] addr_selector2_168;
wire[15:0] addr_remain2_168;
address_decode_4 decoder_2_168 = address_decode_4(addr_selector1_10[8],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_168,addr_remain2_168);


wire[15:0] addr_selector2_169;
wire[15:0] addr_remain2_169;
address_decode_4 decoder_2_169 = address_decode_4(addr_selector1_10[9],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_169,addr_remain2_169);


wire[15:0] addr_selector2_170;
wire[15:0] addr_remain2_170;
address_decode_4 decoder_2_170 = address_decode_4(addr_selector1_10[10],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_170,addr_remain2_170);


wire[15:0] addr_selector2_171;
wire[15:0] addr_remain2_171;
address_decode_4 decoder_2_171 = address_decode_4(addr_selector1_10[11],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_171,addr_remain2_171);


wire[15:0] addr_selector2_172;
wire[15:0] addr_remain2_172;
address_decode_4 decoder_2_172 = address_decode_4(addr_selector1_10[12],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_172,addr_remain2_172);


wire[15:0] addr_selector2_173;
wire[15:0] addr_remain2_173;
address_decode_4 decoder_2_173 = address_decode_4(addr_selector1_10[13],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_173,addr_remain2_173);


wire[15:0] addr_selector2_174;
wire[15:0] addr_remain2_174;
address_decode_4 decoder_2_174 = address_decode_4(addr_selector1_10[14],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_174,addr_remain2_174);


wire[15:0] addr_selector2_175;
wire[15:0] addr_remain2_175;
address_decode_4 decoder_2_175 = address_decode_4(addr_selector1_10[15],addr_remain1_10[31:16],addr_remain1_10,addr_selector2_175,addr_remain2_175);


wire[15:0] addr_selector2_176;
wire[15:0] addr_remain2_176;
address_decode_4 decoder_2_176 = address_decode_4(addr_selector1_11[0],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_176,addr_remain2_176);


wire[15:0] addr_selector2_177;
wire[15:0] addr_remain2_177;
address_decode_4 decoder_2_177 = address_decode_4(addr_selector1_11[1],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_177,addr_remain2_177);


wire[15:0] addr_selector2_178;
wire[15:0] addr_remain2_178;
address_decode_4 decoder_2_178 = address_decode_4(addr_selector1_11[2],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_178,addr_remain2_178);


wire[15:0] addr_selector2_179;
wire[15:0] addr_remain2_179;
address_decode_4 decoder_2_179 = address_decode_4(addr_selector1_11[3],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_179,addr_remain2_179);


wire[15:0] addr_selector2_180;
wire[15:0] addr_remain2_180;
address_decode_4 decoder_2_180 = address_decode_4(addr_selector1_11[4],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_180,addr_remain2_180);


wire[15:0] addr_selector2_181;
wire[15:0] addr_remain2_181;
address_decode_4 decoder_2_181 = address_decode_4(addr_selector1_11[5],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_181,addr_remain2_181);


wire[15:0] addr_selector2_182;
wire[15:0] addr_remain2_182;
address_decode_4 decoder_2_182 = address_decode_4(addr_selector1_11[6],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_182,addr_remain2_182);


wire[15:0] addr_selector2_183;
wire[15:0] addr_remain2_183;
address_decode_4 decoder_2_183 = address_decode_4(addr_selector1_11[7],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_183,addr_remain2_183);


wire[15:0] addr_selector2_184;
wire[15:0] addr_remain2_184;
address_decode_4 decoder_2_184 = address_decode_4(addr_selector1_11[8],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_184,addr_remain2_184);


wire[15:0] addr_selector2_185;
wire[15:0] addr_remain2_185;
address_decode_4 decoder_2_185 = address_decode_4(addr_selector1_11[9],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_185,addr_remain2_185);


wire[15:0] addr_selector2_186;
wire[15:0] addr_remain2_186;
address_decode_4 decoder_2_186 = address_decode_4(addr_selector1_11[10],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_186,addr_remain2_186);


wire[15:0] addr_selector2_187;
wire[15:0] addr_remain2_187;
address_decode_4 decoder_2_187 = address_decode_4(addr_selector1_11[11],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_187,addr_remain2_187);


wire[15:0] addr_selector2_188;
wire[15:0] addr_remain2_188;
address_decode_4 decoder_2_188 = address_decode_4(addr_selector1_11[12],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_188,addr_remain2_188);


wire[15:0] addr_selector2_189;
wire[15:0] addr_remain2_189;
address_decode_4 decoder_2_189 = address_decode_4(addr_selector1_11[13],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_189,addr_remain2_189);


wire[15:0] addr_selector2_190;
wire[15:0] addr_remain2_190;
address_decode_4 decoder_2_190 = address_decode_4(addr_selector1_11[14],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_190,addr_remain2_190);


wire[15:0] addr_selector2_191;
wire[15:0] addr_remain2_191;
address_decode_4 decoder_2_191 = address_decode_4(addr_selector1_11[15],addr_remain1_11[31:16],addr_remain1_11,addr_selector2_191,addr_remain2_191);


wire[15:0] addr_selector2_192;
wire[15:0] addr_remain2_192;
address_decode_4 decoder_2_192 = address_decode_4(addr_selector1_12[0],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_192,addr_remain2_192);


wire[15:0] addr_selector2_193;
wire[15:0] addr_remain2_193;
address_decode_4 decoder_2_193 = address_decode_4(addr_selector1_12[1],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_193,addr_remain2_193);


wire[15:0] addr_selector2_194;
wire[15:0] addr_remain2_194;
address_decode_4 decoder_2_194 = address_decode_4(addr_selector1_12[2],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_194,addr_remain2_194);


wire[15:0] addr_selector2_195;
wire[15:0] addr_remain2_195;
address_decode_4 decoder_2_195 = address_decode_4(addr_selector1_12[3],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_195,addr_remain2_195);


wire[15:0] addr_selector2_196;
wire[15:0] addr_remain2_196;
address_decode_4 decoder_2_196 = address_decode_4(addr_selector1_12[4],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_196,addr_remain2_196);


wire[15:0] addr_selector2_197;
wire[15:0] addr_remain2_197;
address_decode_4 decoder_2_197 = address_decode_4(addr_selector1_12[5],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_197,addr_remain2_197);


wire[15:0] addr_selector2_198;
wire[15:0] addr_remain2_198;
address_decode_4 decoder_2_198 = address_decode_4(addr_selector1_12[6],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_198,addr_remain2_198);


wire[15:0] addr_selector2_199;
wire[15:0] addr_remain2_199;
address_decode_4 decoder_2_199 = address_decode_4(addr_selector1_12[7],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_199,addr_remain2_199);


wire[15:0] addr_selector2_200;
wire[15:0] addr_remain2_200;
address_decode_4 decoder_2_200 = address_decode_4(addr_selector1_12[8],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_200,addr_remain2_200);


wire[15:0] addr_selector2_201;
wire[15:0] addr_remain2_201;
address_decode_4 decoder_2_201 = address_decode_4(addr_selector1_12[9],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_201,addr_remain2_201);


wire[15:0] addr_selector2_202;
wire[15:0] addr_remain2_202;
address_decode_4 decoder_2_202 = address_decode_4(addr_selector1_12[10],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_202,addr_remain2_202);


wire[15:0] addr_selector2_203;
wire[15:0] addr_remain2_203;
address_decode_4 decoder_2_203 = address_decode_4(addr_selector1_12[11],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_203,addr_remain2_203);


wire[15:0] addr_selector2_204;
wire[15:0] addr_remain2_204;
address_decode_4 decoder_2_204 = address_decode_4(addr_selector1_12[12],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_204,addr_remain2_204);


wire[15:0] addr_selector2_205;
wire[15:0] addr_remain2_205;
address_decode_4 decoder_2_205 = address_decode_4(addr_selector1_12[13],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_205,addr_remain2_205);


wire[15:0] addr_selector2_206;
wire[15:0] addr_remain2_206;
address_decode_4 decoder_2_206 = address_decode_4(addr_selector1_12[14],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_206,addr_remain2_206);


wire[15:0] addr_selector2_207;
wire[15:0] addr_remain2_207;
address_decode_4 decoder_2_207 = address_decode_4(addr_selector1_12[15],addr_remain1_12[31:16],addr_remain1_12,addr_selector2_207,addr_remain2_207);


wire[15:0] addr_selector2_208;
wire[15:0] addr_remain2_208;
address_decode_4 decoder_2_208 = address_decode_4(addr_selector1_13[0],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_208,addr_remain2_208);


wire[15:0] addr_selector2_209;
wire[15:0] addr_remain2_209;
address_decode_4 decoder_2_209 = address_decode_4(addr_selector1_13[1],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_209,addr_remain2_209);


wire[15:0] addr_selector2_210;
wire[15:0] addr_remain2_210;
address_decode_4 decoder_2_210 = address_decode_4(addr_selector1_13[2],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_210,addr_remain2_210);


wire[15:0] addr_selector2_211;
wire[15:0] addr_remain2_211;
address_decode_4 decoder_2_211 = address_decode_4(addr_selector1_13[3],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_211,addr_remain2_211);


wire[15:0] addr_selector2_212;
wire[15:0] addr_remain2_212;
address_decode_4 decoder_2_212 = address_decode_4(addr_selector1_13[4],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_212,addr_remain2_212);


wire[15:0] addr_selector2_213;
wire[15:0] addr_remain2_213;
address_decode_4 decoder_2_213 = address_decode_4(addr_selector1_13[5],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_213,addr_remain2_213);


wire[15:0] addr_selector2_214;
wire[15:0] addr_remain2_214;
address_decode_4 decoder_2_214 = address_decode_4(addr_selector1_13[6],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_214,addr_remain2_214);


wire[15:0] addr_selector2_215;
wire[15:0] addr_remain2_215;
address_decode_4 decoder_2_215 = address_decode_4(addr_selector1_13[7],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_215,addr_remain2_215);


wire[15:0] addr_selector2_216;
wire[15:0] addr_remain2_216;
address_decode_4 decoder_2_216 = address_decode_4(addr_selector1_13[8],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_216,addr_remain2_216);


wire[15:0] addr_selector2_217;
wire[15:0] addr_remain2_217;
address_decode_4 decoder_2_217 = address_decode_4(addr_selector1_13[9],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_217,addr_remain2_217);


wire[15:0] addr_selector2_218;
wire[15:0] addr_remain2_218;
address_decode_4 decoder_2_218 = address_decode_4(addr_selector1_13[10],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_218,addr_remain2_218);


wire[15:0] addr_selector2_219;
wire[15:0] addr_remain2_219;
address_decode_4 decoder_2_219 = address_decode_4(addr_selector1_13[11],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_219,addr_remain2_219);


wire[15:0] addr_selector2_220;
wire[15:0] addr_remain2_220;
address_decode_4 decoder_2_220 = address_decode_4(addr_selector1_13[12],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_220,addr_remain2_220);


wire[15:0] addr_selector2_221;
wire[15:0] addr_remain2_221;
address_decode_4 decoder_2_221 = address_decode_4(addr_selector1_13[13],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_221,addr_remain2_221);


wire[15:0] addr_selector2_222;
wire[15:0] addr_remain2_222;
address_decode_4 decoder_2_222 = address_decode_4(addr_selector1_13[14],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_222,addr_remain2_222);


wire[15:0] addr_selector2_223;
wire[15:0] addr_remain2_223;
address_decode_4 decoder_2_223 = address_decode_4(addr_selector1_13[15],addr_remain1_13[31:16],addr_remain1_13,addr_selector2_223,addr_remain2_223);


wire[15:0] addr_selector2_224;
wire[15:0] addr_remain2_224;
address_decode_4 decoder_2_224 = address_decode_4(addr_selector1_14[0],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_224,addr_remain2_224);


wire[15:0] addr_selector2_225;
wire[15:0] addr_remain2_225;
address_decode_4 decoder_2_225 = address_decode_4(addr_selector1_14[1],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_225,addr_remain2_225);


wire[15:0] addr_selector2_226;
wire[15:0] addr_remain2_226;
address_decode_4 decoder_2_226 = address_decode_4(addr_selector1_14[2],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_226,addr_remain2_226);


wire[15:0] addr_selector2_227;
wire[15:0] addr_remain2_227;
address_decode_4 decoder_2_227 = address_decode_4(addr_selector1_14[3],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_227,addr_remain2_227);


wire[15:0] addr_selector2_228;
wire[15:0] addr_remain2_228;
address_decode_4 decoder_2_228 = address_decode_4(addr_selector1_14[4],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_228,addr_remain2_228);


wire[15:0] addr_selector2_229;
wire[15:0] addr_remain2_229;
address_decode_4 decoder_2_229 = address_decode_4(addr_selector1_14[5],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_229,addr_remain2_229);


wire[15:0] addr_selector2_230;
wire[15:0] addr_remain2_230;
address_decode_4 decoder_2_230 = address_decode_4(addr_selector1_14[6],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_230,addr_remain2_230);


wire[15:0] addr_selector2_231;
wire[15:0] addr_remain2_231;
address_decode_4 decoder_2_231 = address_decode_4(addr_selector1_14[7],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_231,addr_remain2_231);


wire[15:0] addr_selector2_232;
wire[15:0] addr_remain2_232;
address_decode_4 decoder_2_232 = address_decode_4(addr_selector1_14[8],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_232,addr_remain2_232);


wire[15:0] addr_selector2_233;
wire[15:0] addr_remain2_233;
address_decode_4 decoder_2_233 = address_decode_4(addr_selector1_14[9],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_233,addr_remain2_233);


wire[15:0] addr_selector2_234;
wire[15:0] addr_remain2_234;
address_decode_4 decoder_2_234 = address_decode_4(addr_selector1_14[10],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_234,addr_remain2_234);


wire[15:0] addr_selector2_235;
wire[15:0] addr_remain2_235;
address_decode_4 decoder_2_235 = address_decode_4(addr_selector1_14[11],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_235,addr_remain2_235);


wire[15:0] addr_selector2_236;
wire[15:0] addr_remain2_236;
address_decode_4 decoder_2_236 = address_decode_4(addr_selector1_14[12],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_236,addr_remain2_236);


wire[15:0] addr_selector2_237;
wire[15:0] addr_remain2_237;
address_decode_4 decoder_2_237 = address_decode_4(addr_selector1_14[13],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_237,addr_remain2_237);


wire[15:0] addr_selector2_238;
wire[15:0] addr_remain2_238;
address_decode_4 decoder_2_238 = address_decode_4(addr_selector1_14[14],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_238,addr_remain2_238);


wire[15:0] addr_selector2_239;
wire[15:0] addr_remain2_239;
address_decode_4 decoder_2_239 = address_decode_4(addr_selector1_14[15],addr_remain1_14[31:16],addr_remain1_14,addr_selector2_239,addr_remain2_239);


wire[15:0] addr_selector2_240;
wire[15:0] addr_remain2_240;
address_decode_4 decoder_2_240 = address_decode_4(addr_selector1_15[0],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_240,addr_remain2_240);


wire[15:0] addr_selector2_241;
wire[15:0] addr_remain2_241;
address_decode_4 decoder_2_241 = address_decode_4(addr_selector1_15[1],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_241,addr_remain2_241);


wire[15:0] addr_selector2_242;
wire[15:0] addr_remain2_242;
address_decode_4 decoder_2_242 = address_decode_4(addr_selector1_15[2],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_242,addr_remain2_242);


wire[15:0] addr_selector2_243;
wire[15:0] addr_remain2_243;
address_decode_4 decoder_2_243 = address_decode_4(addr_selector1_15[3],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_243,addr_remain2_243);


wire[15:0] addr_selector2_244;
wire[15:0] addr_remain2_244;
address_decode_4 decoder_2_244 = address_decode_4(addr_selector1_15[4],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_244,addr_remain2_244);


wire[15:0] addr_selector2_245;
wire[15:0] addr_remain2_245;
address_decode_4 decoder_2_245 = address_decode_4(addr_selector1_15[5],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_245,addr_remain2_245);


wire[15:0] addr_selector2_246;
wire[15:0] addr_remain2_246;
address_decode_4 decoder_2_246 = address_decode_4(addr_selector1_15[6],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_246,addr_remain2_246);


wire[15:0] addr_selector2_247;
wire[15:0] addr_remain2_247;
address_decode_4 decoder_2_247 = address_decode_4(addr_selector1_15[7],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_247,addr_remain2_247);


wire[15:0] addr_selector2_248;
wire[15:0] addr_remain2_248;
address_decode_4 decoder_2_248 = address_decode_4(addr_selector1_15[8],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_248,addr_remain2_248);


wire[15:0] addr_selector2_249;
wire[15:0] addr_remain2_249;
address_decode_4 decoder_2_249 = address_decode_4(addr_selector1_15[9],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_249,addr_remain2_249);


wire[15:0] addr_selector2_250;
wire[15:0] addr_remain2_250;
address_decode_4 decoder_2_250 = address_decode_4(addr_selector1_15[10],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_250,addr_remain2_250);


wire[15:0] addr_selector2_251;
wire[15:0] addr_remain2_251;
address_decode_4 decoder_2_251 = address_decode_4(addr_selector1_15[11],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_251,addr_remain2_251);


wire[15:0] addr_selector2_252;
wire[15:0] addr_remain2_252;
address_decode_4 decoder_2_252 = address_decode_4(addr_selector1_15[12],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_252,addr_remain2_252);


wire[15:0] addr_selector2_253;
wire[15:0] addr_remain2_253;
address_decode_4 decoder_2_253 = address_decode_4(addr_selector1_15[13],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_253,addr_remain2_253);


wire[15:0] addr_selector2_254;
wire[15:0] addr_remain2_254;
address_decode_4 decoder_2_254 = address_decode_4(addr_selector1_15[14],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_254,addr_remain2_254);


wire[15:0] addr_selector2_255;
wire[15:0] addr_remain2_255;
address_decode_4 decoder_2_255 = address_decode_4(addr_selector1_15[15],addr_remain1_15[31:16],addr_remain1_15,addr_selector2_255,addr_remain2_255);


wire[15:0] addr_selector3_0;
wire[15:0] addr_remain3_0;
address_decode_4 decoder_3_0 = address_decode_4(addr_selector2_0[0],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_0,addr_remain3_0);


wire[15:0] addr_selector3_1;
wire[15:0] addr_remain3_1;
address_decode_4 decoder_3_1 = address_decode_4(addr_selector2_0[1],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_1,addr_remain3_1);


wire[15:0] addr_selector3_2;
wire[15:0] addr_remain3_2;
address_decode_4 decoder_3_2 = address_decode_4(addr_selector2_0[2],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_2,addr_remain3_2);


wire[15:0] addr_selector3_3;
wire[15:0] addr_remain3_3;
address_decode_4 decoder_3_3 = address_decode_4(addr_selector2_0[3],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_3,addr_remain3_3);


wire[15:0] addr_selector3_4;
wire[15:0] addr_remain3_4;
address_decode_4 decoder_3_4 = address_decode_4(addr_selector2_0[4],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_4,addr_remain3_4);


wire[15:0] addr_selector3_5;
wire[15:0] addr_remain3_5;
address_decode_4 decoder_3_5 = address_decode_4(addr_selector2_0[5],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_5,addr_remain3_5);


wire[15:0] addr_selector3_6;
wire[15:0] addr_remain3_6;
address_decode_4 decoder_3_6 = address_decode_4(addr_selector2_0[6],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_6,addr_remain3_6);


wire[15:0] addr_selector3_7;
wire[15:0] addr_remain3_7;
address_decode_4 decoder_3_7 = address_decode_4(addr_selector2_0[7],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_7,addr_remain3_7);


wire[15:0] addr_selector3_8;
wire[15:0] addr_remain3_8;
address_decode_4 decoder_3_8 = address_decode_4(addr_selector2_0[8],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_8,addr_remain3_8);


wire[15:0] addr_selector3_9;
wire[15:0] addr_remain3_9;
address_decode_4 decoder_3_9 = address_decode_4(addr_selector2_0[9],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_9,addr_remain3_9);


wire[15:0] addr_selector3_10;
wire[15:0] addr_remain3_10;
address_decode_4 decoder_3_10 = address_decode_4(addr_selector2_0[10],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_10,addr_remain3_10);


wire[15:0] addr_selector3_11;
wire[15:0] addr_remain3_11;
address_decode_4 decoder_3_11 = address_decode_4(addr_selector2_0[11],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_11,addr_remain3_11);


wire[15:0] addr_selector3_12;
wire[15:0] addr_remain3_12;
address_decode_4 decoder_3_12 = address_decode_4(addr_selector2_0[12],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_12,addr_remain3_12);


wire[15:0] addr_selector3_13;
wire[15:0] addr_remain3_13;
address_decode_4 decoder_3_13 = address_decode_4(addr_selector2_0[13],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_13,addr_remain3_13);


wire[15:0] addr_selector3_14;
wire[15:0] addr_remain3_14;
address_decode_4 decoder_3_14 = address_decode_4(addr_selector2_0[14],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_14,addr_remain3_14);


wire[15:0] addr_selector3_15;
wire[15:0] addr_remain3_15;
address_decode_4 decoder_3_15 = address_decode_4(addr_selector2_0[15],addr_remain2_0[15:0],addr_remain2_0,addr_selector3_15,addr_remain3_15);


wire[15:0] addr_selector3_16;
wire[15:0] addr_remain3_16;
address_decode_4 decoder_3_16 = address_decode_4(addr_selector2_1[0],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_16,addr_remain3_16);


wire[15:0] addr_selector3_17;
wire[15:0] addr_remain3_17;
address_decode_4 decoder_3_17 = address_decode_4(addr_selector2_1[1],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_17,addr_remain3_17);


wire[15:0] addr_selector3_18;
wire[15:0] addr_remain3_18;
address_decode_4 decoder_3_18 = address_decode_4(addr_selector2_1[2],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_18,addr_remain3_18);


wire[15:0] addr_selector3_19;
wire[15:0] addr_remain3_19;
address_decode_4 decoder_3_19 = address_decode_4(addr_selector2_1[3],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_19,addr_remain3_19);


wire[15:0] addr_selector3_20;
wire[15:0] addr_remain3_20;
address_decode_4 decoder_3_20 = address_decode_4(addr_selector2_1[4],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_20,addr_remain3_20);


wire[15:0] addr_selector3_21;
wire[15:0] addr_remain3_21;
address_decode_4 decoder_3_21 = address_decode_4(addr_selector2_1[5],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_21,addr_remain3_21);


wire[15:0] addr_selector3_22;
wire[15:0] addr_remain3_22;
address_decode_4 decoder_3_22 = address_decode_4(addr_selector2_1[6],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_22,addr_remain3_22);


wire[15:0] addr_selector3_23;
wire[15:0] addr_remain3_23;
address_decode_4 decoder_3_23 = address_decode_4(addr_selector2_1[7],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_23,addr_remain3_23);


wire[15:0] addr_selector3_24;
wire[15:0] addr_remain3_24;
address_decode_4 decoder_3_24 = address_decode_4(addr_selector2_1[8],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_24,addr_remain3_24);


wire[15:0] addr_selector3_25;
wire[15:0] addr_remain3_25;
address_decode_4 decoder_3_25 = address_decode_4(addr_selector2_1[9],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_25,addr_remain3_25);


wire[15:0] addr_selector3_26;
wire[15:0] addr_remain3_26;
address_decode_4 decoder_3_26 = address_decode_4(addr_selector2_1[10],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_26,addr_remain3_26);


wire[15:0] addr_selector3_27;
wire[15:0] addr_remain3_27;
address_decode_4 decoder_3_27 = address_decode_4(addr_selector2_1[11],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_27,addr_remain3_27);


wire[15:0] addr_selector3_28;
wire[15:0] addr_remain3_28;
address_decode_4 decoder_3_28 = address_decode_4(addr_selector2_1[12],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_28,addr_remain3_28);


wire[15:0] addr_selector3_29;
wire[15:0] addr_remain3_29;
address_decode_4 decoder_3_29 = address_decode_4(addr_selector2_1[13],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_29,addr_remain3_29);


wire[15:0] addr_selector3_30;
wire[15:0] addr_remain3_30;
address_decode_4 decoder_3_30 = address_decode_4(addr_selector2_1[14],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_30,addr_remain3_30);


wire[15:0] addr_selector3_31;
wire[15:0] addr_remain3_31;
address_decode_4 decoder_3_31 = address_decode_4(addr_selector2_1[15],addr_remain2_1[15:0],addr_remain2_1,addr_selector3_31,addr_remain3_31);


wire[15:0] addr_selector3_32;
wire[15:0] addr_remain3_32;
address_decode_4 decoder_3_32 = address_decode_4(addr_selector2_2[0],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_32,addr_remain3_32);


wire[15:0] addr_selector3_33;
wire[15:0] addr_remain3_33;
address_decode_4 decoder_3_33 = address_decode_4(addr_selector2_2[1],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_33,addr_remain3_33);


wire[15:0] addr_selector3_34;
wire[15:0] addr_remain3_34;
address_decode_4 decoder_3_34 = address_decode_4(addr_selector2_2[2],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_34,addr_remain3_34);


wire[15:0] addr_selector3_35;
wire[15:0] addr_remain3_35;
address_decode_4 decoder_3_35 = address_decode_4(addr_selector2_2[3],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_35,addr_remain3_35);


wire[15:0] addr_selector3_36;
wire[15:0] addr_remain3_36;
address_decode_4 decoder_3_36 = address_decode_4(addr_selector2_2[4],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_36,addr_remain3_36);


wire[15:0] addr_selector3_37;
wire[15:0] addr_remain3_37;
address_decode_4 decoder_3_37 = address_decode_4(addr_selector2_2[5],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_37,addr_remain3_37);


wire[15:0] addr_selector3_38;
wire[15:0] addr_remain3_38;
address_decode_4 decoder_3_38 = address_decode_4(addr_selector2_2[6],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_38,addr_remain3_38);


wire[15:0] addr_selector3_39;
wire[15:0] addr_remain3_39;
address_decode_4 decoder_3_39 = address_decode_4(addr_selector2_2[7],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_39,addr_remain3_39);


wire[15:0] addr_selector3_40;
wire[15:0] addr_remain3_40;
address_decode_4 decoder_3_40 = address_decode_4(addr_selector2_2[8],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_40,addr_remain3_40);


wire[15:0] addr_selector3_41;
wire[15:0] addr_remain3_41;
address_decode_4 decoder_3_41 = address_decode_4(addr_selector2_2[9],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_41,addr_remain3_41);


wire[15:0] addr_selector3_42;
wire[15:0] addr_remain3_42;
address_decode_4 decoder_3_42 = address_decode_4(addr_selector2_2[10],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_42,addr_remain3_42);


wire[15:0] addr_selector3_43;
wire[15:0] addr_remain3_43;
address_decode_4 decoder_3_43 = address_decode_4(addr_selector2_2[11],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_43,addr_remain3_43);


wire[15:0] addr_selector3_44;
wire[15:0] addr_remain3_44;
address_decode_4 decoder_3_44 = address_decode_4(addr_selector2_2[12],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_44,addr_remain3_44);


wire[15:0] addr_selector3_45;
wire[15:0] addr_remain3_45;
address_decode_4 decoder_3_45 = address_decode_4(addr_selector2_2[13],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_45,addr_remain3_45);


wire[15:0] addr_selector3_46;
wire[15:0] addr_remain3_46;
address_decode_4 decoder_3_46 = address_decode_4(addr_selector2_2[14],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_46,addr_remain3_46);


wire[15:0] addr_selector3_47;
wire[15:0] addr_remain3_47;
address_decode_4 decoder_3_47 = address_decode_4(addr_selector2_2[15],addr_remain2_2[15:0],addr_remain2_2,addr_selector3_47,addr_remain3_47);


wire[15:0] addr_selector3_48;
wire[15:0] addr_remain3_48;
address_decode_4 decoder_3_48 = address_decode_4(addr_selector2_3[0],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_48,addr_remain3_48);


wire[15:0] addr_selector3_49;
wire[15:0] addr_remain3_49;
address_decode_4 decoder_3_49 = address_decode_4(addr_selector2_3[1],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_49,addr_remain3_49);


wire[15:0] addr_selector3_50;
wire[15:0] addr_remain3_50;
address_decode_4 decoder_3_50 = address_decode_4(addr_selector2_3[2],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_50,addr_remain3_50);


wire[15:0] addr_selector3_51;
wire[15:0] addr_remain3_51;
address_decode_4 decoder_3_51 = address_decode_4(addr_selector2_3[3],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_51,addr_remain3_51);


wire[15:0] addr_selector3_52;
wire[15:0] addr_remain3_52;
address_decode_4 decoder_3_52 = address_decode_4(addr_selector2_3[4],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_52,addr_remain3_52);


wire[15:0] addr_selector3_53;
wire[15:0] addr_remain3_53;
address_decode_4 decoder_3_53 = address_decode_4(addr_selector2_3[5],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_53,addr_remain3_53);


wire[15:0] addr_selector3_54;
wire[15:0] addr_remain3_54;
address_decode_4 decoder_3_54 = address_decode_4(addr_selector2_3[6],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_54,addr_remain3_54);


wire[15:0] addr_selector3_55;
wire[15:0] addr_remain3_55;
address_decode_4 decoder_3_55 = address_decode_4(addr_selector2_3[7],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_55,addr_remain3_55);


wire[15:0] addr_selector3_56;
wire[15:0] addr_remain3_56;
address_decode_4 decoder_3_56 = address_decode_4(addr_selector2_3[8],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_56,addr_remain3_56);


wire[15:0] addr_selector3_57;
wire[15:0] addr_remain3_57;
address_decode_4 decoder_3_57 = address_decode_4(addr_selector2_3[9],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_57,addr_remain3_57);


wire[15:0] addr_selector3_58;
wire[15:0] addr_remain3_58;
address_decode_4 decoder_3_58 = address_decode_4(addr_selector2_3[10],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_58,addr_remain3_58);


wire[15:0] addr_selector3_59;
wire[15:0] addr_remain3_59;
address_decode_4 decoder_3_59 = address_decode_4(addr_selector2_3[11],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_59,addr_remain3_59);


wire[15:0] addr_selector3_60;
wire[15:0] addr_remain3_60;
address_decode_4 decoder_3_60 = address_decode_4(addr_selector2_3[12],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_60,addr_remain3_60);


wire[15:0] addr_selector3_61;
wire[15:0] addr_remain3_61;
address_decode_4 decoder_3_61 = address_decode_4(addr_selector2_3[13],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_61,addr_remain3_61);


wire[15:0] addr_selector3_62;
wire[15:0] addr_remain3_62;
address_decode_4 decoder_3_62 = address_decode_4(addr_selector2_3[14],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_62,addr_remain3_62);


wire[15:0] addr_selector3_63;
wire[15:0] addr_remain3_63;
address_decode_4 decoder_3_63 = address_decode_4(addr_selector2_3[15],addr_remain2_3[15:0],addr_remain2_3,addr_selector3_63,addr_remain3_63);


wire[15:0] addr_selector3_64;
wire[15:0] addr_remain3_64;
address_decode_4 decoder_3_64 = address_decode_4(addr_selector2_4[0],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_64,addr_remain3_64);


wire[15:0] addr_selector3_65;
wire[15:0] addr_remain3_65;
address_decode_4 decoder_3_65 = address_decode_4(addr_selector2_4[1],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_65,addr_remain3_65);


wire[15:0] addr_selector3_66;
wire[15:0] addr_remain3_66;
address_decode_4 decoder_3_66 = address_decode_4(addr_selector2_4[2],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_66,addr_remain3_66);


wire[15:0] addr_selector3_67;
wire[15:0] addr_remain3_67;
address_decode_4 decoder_3_67 = address_decode_4(addr_selector2_4[3],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_67,addr_remain3_67);


wire[15:0] addr_selector3_68;
wire[15:0] addr_remain3_68;
address_decode_4 decoder_3_68 = address_decode_4(addr_selector2_4[4],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_68,addr_remain3_68);


wire[15:0] addr_selector3_69;
wire[15:0] addr_remain3_69;
address_decode_4 decoder_3_69 = address_decode_4(addr_selector2_4[5],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_69,addr_remain3_69);


wire[15:0] addr_selector3_70;
wire[15:0] addr_remain3_70;
address_decode_4 decoder_3_70 = address_decode_4(addr_selector2_4[6],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_70,addr_remain3_70);


wire[15:0] addr_selector3_71;
wire[15:0] addr_remain3_71;
address_decode_4 decoder_3_71 = address_decode_4(addr_selector2_4[7],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_71,addr_remain3_71);


wire[15:0] addr_selector3_72;
wire[15:0] addr_remain3_72;
address_decode_4 decoder_3_72 = address_decode_4(addr_selector2_4[8],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_72,addr_remain3_72);


wire[15:0] addr_selector3_73;
wire[15:0] addr_remain3_73;
address_decode_4 decoder_3_73 = address_decode_4(addr_selector2_4[9],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_73,addr_remain3_73);


wire[15:0] addr_selector3_74;
wire[15:0] addr_remain3_74;
address_decode_4 decoder_3_74 = address_decode_4(addr_selector2_4[10],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_74,addr_remain3_74);


wire[15:0] addr_selector3_75;
wire[15:0] addr_remain3_75;
address_decode_4 decoder_3_75 = address_decode_4(addr_selector2_4[11],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_75,addr_remain3_75);


wire[15:0] addr_selector3_76;
wire[15:0] addr_remain3_76;
address_decode_4 decoder_3_76 = address_decode_4(addr_selector2_4[12],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_76,addr_remain3_76);


wire[15:0] addr_selector3_77;
wire[15:0] addr_remain3_77;
address_decode_4 decoder_3_77 = address_decode_4(addr_selector2_4[13],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_77,addr_remain3_77);


wire[15:0] addr_selector3_78;
wire[15:0] addr_remain3_78;
address_decode_4 decoder_3_78 = address_decode_4(addr_selector2_4[14],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_78,addr_remain3_78);


wire[15:0] addr_selector3_79;
wire[15:0] addr_remain3_79;
address_decode_4 decoder_3_79 = address_decode_4(addr_selector2_4[15],addr_remain2_4[15:0],addr_remain2_4,addr_selector3_79,addr_remain3_79);


wire[15:0] addr_selector3_80;
wire[15:0] addr_remain3_80;
address_decode_4 decoder_3_80 = address_decode_4(addr_selector2_5[0],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_80,addr_remain3_80);


wire[15:0] addr_selector3_81;
wire[15:0] addr_remain3_81;
address_decode_4 decoder_3_81 = address_decode_4(addr_selector2_5[1],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_81,addr_remain3_81);


wire[15:0] addr_selector3_82;
wire[15:0] addr_remain3_82;
address_decode_4 decoder_3_82 = address_decode_4(addr_selector2_5[2],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_82,addr_remain3_82);


wire[15:0] addr_selector3_83;
wire[15:0] addr_remain3_83;
address_decode_4 decoder_3_83 = address_decode_4(addr_selector2_5[3],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_83,addr_remain3_83);


wire[15:0] addr_selector3_84;
wire[15:0] addr_remain3_84;
address_decode_4 decoder_3_84 = address_decode_4(addr_selector2_5[4],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_84,addr_remain3_84);


wire[15:0] addr_selector3_85;
wire[15:0] addr_remain3_85;
address_decode_4 decoder_3_85 = address_decode_4(addr_selector2_5[5],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_85,addr_remain3_85);


wire[15:0] addr_selector3_86;
wire[15:0] addr_remain3_86;
address_decode_4 decoder_3_86 = address_decode_4(addr_selector2_5[6],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_86,addr_remain3_86);


wire[15:0] addr_selector3_87;
wire[15:0] addr_remain3_87;
address_decode_4 decoder_3_87 = address_decode_4(addr_selector2_5[7],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_87,addr_remain3_87);


wire[15:0] addr_selector3_88;
wire[15:0] addr_remain3_88;
address_decode_4 decoder_3_88 = address_decode_4(addr_selector2_5[8],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_88,addr_remain3_88);


wire[15:0] addr_selector3_89;
wire[15:0] addr_remain3_89;
address_decode_4 decoder_3_89 = address_decode_4(addr_selector2_5[9],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_89,addr_remain3_89);


wire[15:0] addr_selector3_90;
wire[15:0] addr_remain3_90;
address_decode_4 decoder_3_90 = address_decode_4(addr_selector2_5[10],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_90,addr_remain3_90);


wire[15:0] addr_selector3_91;
wire[15:0] addr_remain3_91;
address_decode_4 decoder_3_91 = address_decode_4(addr_selector2_5[11],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_91,addr_remain3_91);


wire[15:0] addr_selector3_92;
wire[15:0] addr_remain3_92;
address_decode_4 decoder_3_92 = address_decode_4(addr_selector2_5[12],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_92,addr_remain3_92);


wire[15:0] addr_selector3_93;
wire[15:0] addr_remain3_93;
address_decode_4 decoder_3_93 = address_decode_4(addr_selector2_5[13],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_93,addr_remain3_93);


wire[15:0] addr_selector3_94;
wire[15:0] addr_remain3_94;
address_decode_4 decoder_3_94 = address_decode_4(addr_selector2_5[14],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_94,addr_remain3_94);


wire[15:0] addr_selector3_95;
wire[15:0] addr_remain3_95;
address_decode_4 decoder_3_95 = address_decode_4(addr_selector2_5[15],addr_remain2_5[15:0],addr_remain2_5,addr_selector3_95,addr_remain3_95);


wire[15:0] addr_selector3_96;
wire[15:0] addr_remain3_96;
address_decode_4 decoder_3_96 = address_decode_4(addr_selector2_6[0],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_96,addr_remain3_96);


wire[15:0] addr_selector3_97;
wire[15:0] addr_remain3_97;
address_decode_4 decoder_3_97 = address_decode_4(addr_selector2_6[1],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_97,addr_remain3_97);


wire[15:0] addr_selector3_98;
wire[15:0] addr_remain3_98;
address_decode_4 decoder_3_98 = address_decode_4(addr_selector2_6[2],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_98,addr_remain3_98);


wire[15:0] addr_selector3_99;
wire[15:0] addr_remain3_99;
address_decode_4 decoder_3_99 = address_decode_4(addr_selector2_6[3],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_99,addr_remain3_99);


wire[15:0] addr_selector3_100;
wire[15:0] addr_remain3_100;
address_decode_4 decoder_3_100 = address_decode_4(addr_selector2_6[4],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_100,addr_remain3_100);


wire[15:0] addr_selector3_101;
wire[15:0] addr_remain3_101;
address_decode_4 decoder_3_101 = address_decode_4(addr_selector2_6[5],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_101,addr_remain3_101);


wire[15:0] addr_selector3_102;
wire[15:0] addr_remain3_102;
address_decode_4 decoder_3_102 = address_decode_4(addr_selector2_6[6],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_102,addr_remain3_102);


wire[15:0] addr_selector3_103;
wire[15:0] addr_remain3_103;
address_decode_4 decoder_3_103 = address_decode_4(addr_selector2_6[7],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_103,addr_remain3_103);


wire[15:0] addr_selector3_104;
wire[15:0] addr_remain3_104;
address_decode_4 decoder_3_104 = address_decode_4(addr_selector2_6[8],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_104,addr_remain3_104);


wire[15:0] addr_selector3_105;
wire[15:0] addr_remain3_105;
address_decode_4 decoder_3_105 = address_decode_4(addr_selector2_6[9],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_105,addr_remain3_105);


wire[15:0] addr_selector3_106;
wire[15:0] addr_remain3_106;
address_decode_4 decoder_3_106 = address_decode_4(addr_selector2_6[10],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_106,addr_remain3_106);


wire[15:0] addr_selector3_107;
wire[15:0] addr_remain3_107;
address_decode_4 decoder_3_107 = address_decode_4(addr_selector2_6[11],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_107,addr_remain3_107);


wire[15:0] addr_selector3_108;
wire[15:0] addr_remain3_108;
address_decode_4 decoder_3_108 = address_decode_4(addr_selector2_6[12],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_108,addr_remain3_108);


wire[15:0] addr_selector3_109;
wire[15:0] addr_remain3_109;
address_decode_4 decoder_3_109 = address_decode_4(addr_selector2_6[13],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_109,addr_remain3_109);


wire[15:0] addr_selector3_110;
wire[15:0] addr_remain3_110;
address_decode_4 decoder_3_110 = address_decode_4(addr_selector2_6[14],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_110,addr_remain3_110);


wire[15:0] addr_selector3_111;
wire[15:0] addr_remain3_111;
address_decode_4 decoder_3_111 = address_decode_4(addr_selector2_6[15],addr_remain2_6[15:0],addr_remain2_6,addr_selector3_111,addr_remain3_111);


wire[15:0] addr_selector3_112;
wire[15:0] addr_remain3_112;
address_decode_4 decoder_3_112 = address_decode_4(addr_selector2_7[0],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_112,addr_remain3_112);


wire[15:0] addr_selector3_113;
wire[15:0] addr_remain3_113;
address_decode_4 decoder_3_113 = address_decode_4(addr_selector2_7[1],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_113,addr_remain3_113);


wire[15:0] addr_selector3_114;
wire[15:0] addr_remain3_114;
address_decode_4 decoder_3_114 = address_decode_4(addr_selector2_7[2],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_114,addr_remain3_114);


wire[15:0] addr_selector3_115;
wire[15:0] addr_remain3_115;
address_decode_4 decoder_3_115 = address_decode_4(addr_selector2_7[3],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_115,addr_remain3_115);


wire[15:0] addr_selector3_116;
wire[15:0] addr_remain3_116;
address_decode_4 decoder_3_116 = address_decode_4(addr_selector2_7[4],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_116,addr_remain3_116);


wire[15:0] addr_selector3_117;
wire[15:0] addr_remain3_117;
address_decode_4 decoder_3_117 = address_decode_4(addr_selector2_7[5],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_117,addr_remain3_117);


wire[15:0] addr_selector3_118;
wire[15:0] addr_remain3_118;
address_decode_4 decoder_3_118 = address_decode_4(addr_selector2_7[6],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_118,addr_remain3_118);


wire[15:0] addr_selector3_119;
wire[15:0] addr_remain3_119;
address_decode_4 decoder_3_119 = address_decode_4(addr_selector2_7[7],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_119,addr_remain3_119);


wire[15:0] addr_selector3_120;
wire[15:0] addr_remain3_120;
address_decode_4 decoder_3_120 = address_decode_4(addr_selector2_7[8],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_120,addr_remain3_120);


wire[15:0] addr_selector3_121;
wire[15:0] addr_remain3_121;
address_decode_4 decoder_3_121 = address_decode_4(addr_selector2_7[9],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_121,addr_remain3_121);


wire[15:0] addr_selector3_122;
wire[15:0] addr_remain3_122;
address_decode_4 decoder_3_122 = address_decode_4(addr_selector2_7[10],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_122,addr_remain3_122);


wire[15:0] addr_selector3_123;
wire[15:0] addr_remain3_123;
address_decode_4 decoder_3_123 = address_decode_4(addr_selector2_7[11],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_123,addr_remain3_123);


wire[15:0] addr_selector3_124;
wire[15:0] addr_remain3_124;
address_decode_4 decoder_3_124 = address_decode_4(addr_selector2_7[12],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_124,addr_remain3_124);


wire[15:0] addr_selector3_125;
wire[15:0] addr_remain3_125;
address_decode_4 decoder_3_125 = address_decode_4(addr_selector2_7[13],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_125,addr_remain3_125);


wire[15:0] addr_selector3_126;
wire[15:0] addr_remain3_126;
address_decode_4 decoder_3_126 = address_decode_4(addr_selector2_7[14],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_126,addr_remain3_126);


wire[15:0] addr_selector3_127;
wire[15:0] addr_remain3_127;
address_decode_4 decoder_3_127 = address_decode_4(addr_selector2_7[15],addr_remain2_7[15:0],addr_remain2_7,addr_selector3_127,addr_remain3_127);


wire[15:0] addr_selector3_128;
wire[15:0] addr_remain3_128;
address_decode_4 decoder_3_128 = address_decode_4(addr_selector2_8[0],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_128,addr_remain3_128);


wire[15:0] addr_selector3_129;
wire[15:0] addr_remain3_129;
address_decode_4 decoder_3_129 = address_decode_4(addr_selector2_8[1],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_129,addr_remain3_129);


wire[15:0] addr_selector3_130;
wire[15:0] addr_remain3_130;
address_decode_4 decoder_3_130 = address_decode_4(addr_selector2_8[2],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_130,addr_remain3_130);


wire[15:0] addr_selector3_131;
wire[15:0] addr_remain3_131;
address_decode_4 decoder_3_131 = address_decode_4(addr_selector2_8[3],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_131,addr_remain3_131);


wire[15:0] addr_selector3_132;
wire[15:0] addr_remain3_132;
address_decode_4 decoder_3_132 = address_decode_4(addr_selector2_8[4],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_132,addr_remain3_132);


wire[15:0] addr_selector3_133;
wire[15:0] addr_remain3_133;
address_decode_4 decoder_3_133 = address_decode_4(addr_selector2_8[5],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_133,addr_remain3_133);


wire[15:0] addr_selector3_134;
wire[15:0] addr_remain3_134;
address_decode_4 decoder_3_134 = address_decode_4(addr_selector2_8[6],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_134,addr_remain3_134);


wire[15:0] addr_selector3_135;
wire[15:0] addr_remain3_135;
address_decode_4 decoder_3_135 = address_decode_4(addr_selector2_8[7],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_135,addr_remain3_135);


wire[15:0] addr_selector3_136;
wire[15:0] addr_remain3_136;
address_decode_4 decoder_3_136 = address_decode_4(addr_selector2_8[8],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_136,addr_remain3_136);


wire[15:0] addr_selector3_137;
wire[15:0] addr_remain3_137;
address_decode_4 decoder_3_137 = address_decode_4(addr_selector2_8[9],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_137,addr_remain3_137);


wire[15:0] addr_selector3_138;
wire[15:0] addr_remain3_138;
address_decode_4 decoder_3_138 = address_decode_4(addr_selector2_8[10],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_138,addr_remain3_138);


wire[15:0] addr_selector3_139;
wire[15:0] addr_remain3_139;
address_decode_4 decoder_3_139 = address_decode_4(addr_selector2_8[11],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_139,addr_remain3_139);


wire[15:0] addr_selector3_140;
wire[15:0] addr_remain3_140;
address_decode_4 decoder_3_140 = address_decode_4(addr_selector2_8[12],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_140,addr_remain3_140);


wire[15:0] addr_selector3_141;
wire[15:0] addr_remain3_141;
address_decode_4 decoder_3_141 = address_decode_4(addr_selector2_8[13],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_141,addr_remain3_141);


wire[15:0] addr_selector3_142;
wire[15:0] addr_remain3_142;
address_decode_4 decoder_3_142 = address_decode_4(addr_selector2_8[14],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_142,addr_remain3_142);


wire[15:0] addr_selector3_143;
wire[15:0] addr_remain3_143;
address_decode_4 decoder_3_143 = address_decode_4(addr_selector2_8[15],addr_remain2_8[15:0],addr_remain2_8,addr_selector3_143,addr_remain3_143);


wire[15:0] addr_selector3_144;
wire[15:0] addr_remain3_144;
address_decode_4 decoder_3_144 = address_decode_4(addr_selector2_9[0],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_144,addr_remain3_144);


wire[15:0] addr_selector3_145;
wire[15:0] addr_remain3_145;
address_decode_4 decoder_3_145 = address_decode_4(addr_selector2_9[1],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_145,addr_remain3_145);


wire[15:0] addr_selector3_146;
wire[15:0] addr_remain3_146;
address_decode_4 decoder_3_146 = address_decode_4(addr_selector2_9[2],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_146,addr_remain3_146);


wire[15:0] addr_selector3_147;
wire[15:0] addr_remain3_147;
address_decode_4 decoder_3_147 = address_decode_4(addr_selector2_9[3],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_147,addr_remain3_147);


wire[15:0] addr_selector3_148;
wire[15:0] addr_remain3_148;
address_decode_4 decoder_3_148 = address_decode_4(addr_selector2_9[4],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_148,addr_remain3_148);


wire[15:0] addr_selector3_149;
wire[15:0] addr_remain3_149;
address_decode_4 decoder_3_149 = address_decode_4(addr_selector2_9[5],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_149,addr_remain3_149);


wire[15:0] addr_selector3_150;
wire[15:0] addr_remain3_150;
address_decode_4 decoder_3_150 = address_decode_4(addr_selector2_9[6],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_150,addr_remain3_150);


wire[15:0] addr_selector3_151;
wire[15:0] addr_remain3_151;
address_decode_4 decoder_3_151 = address_decode_4(addr_selector2_9[7],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_151,addr_remain3_151);


wire[15:0] addr_selector3_152;
wire[15:0] addr_remain3_152;
address_decode_4 decoder_3_152 = address_decode_4(addr_selector2_9[8],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_152,addr_remain3_152);


wire[15:0] addr_selector3_153;
wire[15:0] addr_remain3_153;
address_decode_4 decoder_3_153 = address_decode_4(addr_selector2_9[9],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_153,addr_remain3_153);


wire[15:0] addr_selector3_154;
wire[15:0] addr_remain3_154;
address_decode_4 decoder_3_154 = address_decode_4(addr_selector2_9[10],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_154,addr_remain3_154);


wire[15:0] addr_selector3_155;
wire[15:0] addr_remain3_155;
address_decode_4 decoder_3_155 = address_decode_4(addr_selector2_9[11],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_155,addr_remain3_155);


wire[15:0] addr_selector3_156;
wire[15:0] addr_remain3_156;
address_decode_4 decoder_3_156 = address_decode_4(addr_selector2_9[12],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_156,addr_remain3_156);


wire[15:0] addr_selector3_157;
wire[15:0] addr_remain3_157;
address_decode_4 decoder_3_157 = address_decode_4(addr_selector2_9[13],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_157,addr_remain3_157);


wire[15:0] addr_selector3_158;
wire[15:0] addr_remain3_158;
address_decode_4 decoder_3_158 = address_decode_4(addr_selector2_9[14],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_158,addr_remain3_158);


wire[15:0] addr_selector3_159;
wire[15:0] addr_remain3_159;
address_decode_4 decoder_3_159 = address_decode_4(addr_selector2_9[15],addr_remain2_9[15:0],addr_remain2_9,addr_selector3_159,addr_remain3_159);


wire[15:0] addr_selector3_160;
wire[15:0] addr_remain3_160;
address_decode_4 decoder_3_160 = address_decode_4(addr_selector2_10[0],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_160,addr_remain3_160);


wire[15:0] addr_selector3_161;
wire[15:0] addr_remain3_161;
address_decode_4 decoder_3_161 = address_decode_4(addr_selector2_10[1],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_161,addr_remain3_161);


wire[15:0] addr_selector3_162;
wire[15:0] addr_remain3_162;
address_decode_4 decoder_3_162 = address_decode_4(addr_selector2_10[2],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_162,addr_remain3_162);


wire[15:0] addr_selector3_163;
wire[15:0] addr_remain3_163;
address_decode_4 decoder_3_163 = address_decode_4(addr_selector2_10[3],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_163,addr_remain3_163);


wire[15:0] addr_selector3_164;
wire[15:0] addr_remain3_164;
address_decode_4 decoder_3_164 = address_decode_4(addr_selector2_10[4],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_164,addr_remain3_164);


wire[15:0] addr_selector3_165;
wire[15:0] addr_remain3_165;
address_decode_4 decoder_3_165 = address_decode_4(addr_selector2_10[5],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_165,addr_remain3_165);


wire[15:0] addr_selector3_166;
wire[15:0] addr_remain3_166;
address_decode_4 decoder_3_166 = address_decode_4(addr_selector2_10[6],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_166,addr_remain3_166);


wire[15:0] addr_selector3_167;
wire[15:0] addr_remain3_167;
address_decode_4 decoder_3_167 = address_decode_4(addr_selector2_10[7],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_167,addr_remain3_167);


wire[15:0] addr_selector3_168;
wire[15:0] addr_remain3_168;
address_decode_4 decoder_3_168 = address_decode_4(addr_selector2_10[8],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_168,addr_remain3_168);


wire[15:0] addr_selector3_169;
wire[15:0] addr_remain3_169;
address_decode_4 decoder_3_169 = address_decode_4(addr_selector2_10[9],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_169,addr_remain3_169);


wire[15:0] addr_selector3_170;
wire[15:0] addr_remain3_170;
address_decode_4 decoder_3_170 = address_decode_4(addr_selector2_10[10],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_170,addr_remain3_170);


wire[15:0] addr_selector3_171;
wire[15:0] addr_remain3_171;
address_decode_4 decoder_3_171 = address_decode_4(addr_selector2_10[11],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_171,addr_remain3_171);


wire[15:0] addr_selector3_172;
wire[15:0] addr_remain3_172;
address_decode_4 decoder_3_172 = address_decode_4(addr_selector2_10[12],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_172,addr_remain3_172);


wire[15:0] addr_selector3_173;
wire[15:0] addr_remain3_173;
address_decode_4 decoder_3_173 = address_decode_4(addr_selector2_10[13],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_173,addr_remain3_173);


wire[15:0] addr_selector3_174;
wire[15:0] addr_remain3_174;
address_decode_4 decoder_3_174 = address_decode_4(addr_selector2_10[14],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_174,addr_remain3_174);


wire[15:0] addr_selector3_175;
wire[15:0] addr_remain3_175;
address_decode_4 decoder_3_175 = address_decode_4(addr_selector2_10[15],addr_remain2_10[15:0],addr_remain2_10,addr_selector3_175,addr_remain3_175);


wire[15:0] addr_selector3_176;
wire[15:0] addr_remain3_176;
address_decode_4 decoder_3_176 = address_decode_4(addr_selector2_11[0],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_176,addr_remain3_176);


wire[15:0] addr_selector3_177;
wire[15:0] addr_remain3_177;
address_decode_4 decoder_3_177 = address_decode_4(addr_selector2_11[1],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_177,addr_remain3_177);


wire[15:0] addr_selector3_178;
wire[15:0] addr_remain3_178;
address_decode_4 decoder_3_178 = address_decode_4(addr_selector2_11[2],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_178,addr_remain3_178);


wire[15:0] addr_selector3_179;
wire[15:0] addr_remain3_179;
address_decode_4 decoder_3_179 = address_decode_4(addr_selector2_11[3],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_179,addr_remain3_179);


wire[15:0] addr_selector3_180;
wire[15:0] addr_remain3_180;
address_decode_4 decoder_3_180 = address_decode_4(addr_selector2_11[4],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_180,addr_remain3_180);


wire[15:0] addr_selector3_181;
wire[15:0] addr_remain3_181;
address_decode_4 decoder_3_181 = address_decode_4(addr_selector2_11[5],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_181,addr_remain3_181);


wire[15:0] addr_selector3_182;
wire[15:0] addr_remain3_182;
address_decode_4 decoder_3_182 = address_decode_4(addr_selector2_11[6],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_182,addr_remain3_182);


wire[15:0] addr_selector3_183;
wire[15:0] addr_remain3_183;
address_decode_4 decoder_3_183 = address_decode_4(addr_selector2_11[7],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_183,addr_remain3_183);


wire[15:0] addr_selector3_184;
wire[15:0] addr_remain3_184;
address_decode_4 decoder_3_184 = address_decode_4(addr_selector2_11[8],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_184,addr_remain3_184);


wire[15:0] addr_selector3_185;
wire[15:0] addr_remain3_185;
address_decode_4 decoder_3_185 = address_decode_4(addr_selector2_11[9],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_185,addr_remain3_185);


wire[15:0] addr_selector3_186;
wire[15:0] addr_remain3_186;
address_decode_4 decoder_3_186 = address_decode_4(addr_selector2_11[10],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_186,addr_remain3_186);


wire[15:0] addr_selector3_187;
wire[15:0] addr_remain3_187;
address_decode_4 decoder_3_187 = address_decode_4(addr_selector2_11[11],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_187,addr_remain3_187);


wire[15:0] addr_selector3_188;
wire[15:0] addr_remain3_188;
address_decode_4 decoder_3_188 = address_decode_4(addr_selector2_11[12],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_188,addr_remain3_188);


wire[15:0] addr_selector3_189;
wire[15:0] addr_remain3_189;
address_decode_4 decoder_3_189 = address_decode_4(addr_selector2_11[13],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_189,addr_remain3_189);


wire[15:0] addr_selector3_190;
wire[15:0] addr_remain3_190;
address_decode_4 decoder_3_190 = address_decode_4(addr_selector2_11[14],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_190,addr_remain3_190);


wire[15:0] addr_selector3_191;
wire[15:0] addr_remain3_191;
address_decode_4 decoder_3_191 = address_decode_4(addr_selector2_11[15],addr_remain2_11[15:0],addr_remain2_11,addr_selector3_191,addr_remain3_191);


wire[15:0] addr_selector3_192;
wire[15:0] addr_remain3_192;
address_decode_4 decoder_3_192 = address_decode_4(addr_selector2_12[0],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_192,addr_remain3_192);


wire[15:0] addr_selector3_193;
wire[15:0] addr_remain3_193;
address_decode_4 decoder_3_193 = address_decode_4(addr_selector2_12[1],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_193,addr_remain3_193);


wire[15:0] addr_selector3_194;
wire[15:0] addr_remain3_194;
address_decode_4 decoder_3_194 = address_decode_4(addr_selector2_12[2],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_194,addr_remain3_194);


wire[15:0] addr_selector3_195;
wire[15:0] addr_remain3_195;
address_decode_4 decoder_3_195 = address_decode_4(addr_selector2_12[3],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_195,addr_remain3_195);


wire[15:0] addr_selector3_196;
wire[15:0] addr_remain3_196;
address_decode_4 decoder_3_196 = address_decode_4(addr_selector2_12[4],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_196,addr_remain3_196);


wire[15:0] addr_selector3_197;
wire[15:0] addr_remain3_197;
address_decode_4 decoder_3_197 = address_decode_4(addr_selector2_12[5],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_197,addr_remain3_197);


wire[15:0] addr_selector3_198;
wire[15:0] addr_remain3_198;
address_decode_4 decoder_3_198 = address_decode_4(addr_selector2_12[6],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_198,addr_remain3_198);


wire[15:0] addr_selector3_199;
wire[15:0] addr_remain3_199;
address_decode_4 decoder_3_199 = address_decode_4(addr_selector2_12[7],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_199,addr_remain3_199);


wire[15:0] addr_selector3_200;
wire[15:0] addr_remain3_200;
address_decode_4 decoder_3_200 = address_decode_4(addr_selector2_12[8],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_200,addr_remain3_200);


wire[15:0] addr_selector3_201;
wire[15:0] addr_remain3_201;
address_decode_4 decoder_3_201 = address_decode_4(addr_selector2_12[9],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_201,addr_remain3_201);


wire[15:0] addr_selector3_202;
wire[15:0] addr_remain3_202;
address_decode_4 decoder_3_202 = address_decode_4(addr_selector2_12[10],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_202,addr_remain3_202);


wire[15:0] addr_selector3_203;
wire[15:0] addr_remain3_203;
address_decode_4 decoder_3_203 = address_decode_4(addr_selector2_12[11],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_203,addr_remain3_203);


wire[15:0] addr_selector3_204;
wire[15:0] addr_remain3_204;
address_decode_4 decoder_3_204 = address_decode_4(addr_selector2_12[12],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_204,addr_remain3_204);


wire[15:0] addr_selector3_205;
wire[15:0] addr_remain3_205;
address_decode_4 decoder_3_205 = address_decode_4(addr_selector2_12[13],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_205,addr_remain3_205);


wire[15:0] addr_selector3_206;
wire[15:0] addr_remain3_206;
address_decode_4 decoder_3_206 = address_decode_4(addr_selector2_12[14],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_206,addr_remain3_206);


wire[15:0] addr_selector3_207;
wire[15:0] addr_remain3_207;
address_decode_4 decoder_3_207 = address_decode_4(addr_selector2_12[15],addr_remain2_12[15:0],addr_remain2_12,addr_selector3_207,addr_remain3_207);


wire[15:0] addr_selector3_208;
wire[15:0] addr_remain3_208;
address_decode_4 decoder_3_208 = address_decode_4(addr_selector2_13[0],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_208,addr_remain3_208);


wire[15:0] addr_selector3_209;
wire[15:0] addr_remain3_209;
address_decode_4 decoder_3_209 = address_decode_4(addr_selector2_13[1],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_209,addr_remain3_209);


wire[15:0] addr_selector3_210;
wire[15:0] addr_remain3_210;
address_decode_4 decoder_3_210 = address_decode_4(addr_selector2_13[2],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_210,addr_remain3_210);


wire[15:0] addr_selector3_211;
wire[15:0] addr_remain3_211;
address_decode_4 decoder_3_211 = address_decode_4(addr_selector2_13[3],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_211,addr_remain3_211);


wire[15:0] addr_selector3_212;
wire[15:0] addr_remain3_212;
address_decode_4 decoder_3_212 = address_decode_4(addr_selector2_13[4],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_212,addr_remain3_212);


wire[15:0] addr_selector3_213;
wire[15:0] addr_remain3_213;
address_decode_4 decoder_3_213 = address_decode_4(addr_selector2_13[5],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_213,addr_remain3_213);


wire[15:0] addr_selector3_214;
wire[15:0] addr_remain3_214;
address_decode_4 decoder_3_214 = address_decode_4(addr_selector2_13[6],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_214,addr_remain3_214);


wire[15:0] addr_selector3_215;
wire[15:0] addr_remain3_215;
address_decode_4 decoder_3_215 = address_decode_4(addr_selector2_13[7],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_215,addr_remain3_215);


wire[15:0] addr_selector3_216;
wire[15:0] addr_remain3_216;
address_decode_4 decoder_3_216 = address_decode_4(addr_selector2_13[8],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_216,addr_remain3_216);


wire[15:0] addr_selector3_217;
wire[15:0] addr_remain3_217;
address_decode_4 decoder_3_217 = address_decode_4(addr_selector2_13[9],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_217,addr_remain3_217);


wire[15:0] addr_selector3_218;
wire[15:0] addr_remain3_218;
address_decode_4 decoder_3_218 = address_decode_4(addr_selector2_13[10],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_218,addr_remain3_218);


wire[15:0] addr_selector3_219;
wire[15:0] addr_remain3_219;
address_decode_4 decoder_3_219 = address_decode_4(addr_selector2_13[11],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_219,addr_remain3_219);


wire[15:0] addr_selector3_220;
wire[15:0] addr_remain3_220;
address_decode_4 decoder_3_220 = address_decode_4(addr_selector2_13[12],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_220,addr_remain3_220);


wire[15:0] addr_selector3_221;
wire[15:0] addr_remain3_221;
address_decode_4 decoder_3_221 = address_decode_4(addr_selector2_13[13],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_221,addr_remain3_221);


wire[15:0] addr_selector3_222;
wire[15:0] addr_remain3_222;
address_decode_4 decoder_3_222 = address_decode_4(addr_selector2_13[14],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_222,addr_remain3_222);


wire[15:0] addr_selector3_223;
wire[15:0] addr_remain3_223;
address_decode_4 decoder_3_223 = address_decode_4(addr_selector2_13[15],addr_remain2_13[15:0],addr_remain2_13,addr_selector3_223,addr_remain3_223);


wire[15:0] addr_selector3_224;
wire[15:0] addr_remain3_224;
address_decode_4 decoder_3_224 = address_decode_4(addr_selector2_14[0],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_224,addr_remain3_224);


wire[15:0] addr_selector3_225;
wire[15:0] addr_remain3_225;
address_decode_4 decoder_3_225 = address_decode_4(addr_selector2_14[1],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_225,addr_remain3_225);


wire[15:0] addr_selector3_226;
wire[15:0] addr_remain3_226;
address_decode_4 decoder_3_226 = address_decode_4(addr_selector2_14[2],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_226,addr_remain3_226);


wire[15:0] addr_selector3_227;
wire[15:0] addr_remain3_227;
address_decode_4 decoder_3_227 = address_decode_4(addr_selector2_14[3],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_227,addr_remain3_227);


wire[15:0] addr_selector3_228;
wire[15:0] addr_remain3_228;
address_decode_4 decoder_3_228 = address_decode_4(addr_selector2_14[4],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_228,addr_remain3_228);


wire[15:0] addr_selector3_229;
wire[15:0] addr_remain3_229;
address_decode_4 decoder_3_229 = address_decode_4(addr_selector2_14[5],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_229,addr_remain3_229);


wire[15:0] addr_selector3_230;
wire[15:0] addr_remain3_230;
address_decode_4 decoder_3_230 = address_decode_4(addr_selector2_14[6],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_230,addr_remain3_230);


wire[15:0] addr_selector3_231;
wire[15:0] addr_remain3_231;
address_decode_4 decoder_3_231 = address_decode_4(addr_selector2_14[7],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_231,addr_remain3_231);


wire[15:0] addr_selector3_232;
wire[15:0] addr_remain3_232;
address_decode_4 decoder_3_232 = address_decode_4(addr_selector2_14[8],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_232,addr_remain3_232);


wire[15:0] addr_selector3_233;
wire[15:0] addr_remain3_233;
address_decode_4 decoder_3_233 = address_decode_4(addr_selector2_14[9],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_233,addr_remain3_233);


wire[15:0] addr_selector3_234;
wire[15:0] addr_remain3_234;
address_decode_4 decoder_3_234 = address_decode_4(addr_selector2_14[10],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_234,addr_remain3_234);


wire[15:0] addr_selector3_235;
wire[15:0] addr_remain3_235;
address_decode_4 decoder_3_235 = address_decode_4(addr_selector2_14[11],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_235,addr_remain3_235);


wire[15:0] addr_selector3_236;
wire[15:0] addr_remain3_236;
address_decode_4 decoder_3_236 = address_decode_4(addr_selector2_14[12],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_236,addr_remain3_236);


wire[15:0] addr_selector3_237;
wire[15:0] addr_remain3_237;
address_decode_4 decoder_3_237 = address_decode_4(addr_selector2_14[13],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_237,addr_remain3_237);


wire[15:0] addr_selector3_238;
wire[15:0] addr_remain3_238;
address_decode_4 decoder_3_238 = address_decode_4(addr_selector2_14[14],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_238,addr_remain3_238);


wire[15:0] addr_selector3_239;
wire[15:0] addr_remain3_239;
address_decode_4 decoder_3_239 = address_decode_4(addr_selector2_14[15],addr_remain2_14[15:0],addr_remain2_14,addr_selector3_239,addr_remain3_239);


wire[15:0] addr_selector3_240;
wire[15:0] addr_remain3_240;
address_decode_4 decoder_3_240 = address_decode_4(addr_selector2_15[0],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_240,addr_remain3_240);


wire[15:0] addr_selector3_241;
wire[15:0] addr_remain3_241;
address_decode_4 decoder_3_241 = address_decode_4(addr_selector2_15[1],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_241,addr_remain3_241);


wire[15:0] addr_selector3_242;
wire[15:0] addr_remain3_242;
address_decode_4 decoder_3_242 = address_decode_4(addr_selector2_15[2],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_242,addr_remain3_242);


wire[15:0] addr_selector3_243;
wire[15:0] addr_remain3_243;
address_decode_4 decoder_3_243 = address_decode_4(addr_selector2_15[3],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_243,addr_remain3_243);


wire[15:0] addr_selector3_244;
wire[15:0] addr_remain3_244;
address_decode_4 decoder_3_244 = address_decode_4(addr_selector2_15[4],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_244,addr_remain3_244);


wire[15:0] addr_selector3_245;
wire[15:0] addr_remain3_245;
address_decode_4 decoder_3_245 = address_decode_4(addr_selector2_15[5],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_245,addr_remain3_245);


wire[15:0] addr_selector3_246;
wire[15:0] addr_remain3_246;
address_decode_4 decoder_3_246 = address_decode_4(addr_selector2_15[6],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_246,addr_remain3_246);


wire[15:0] addr_selector3_247;
wire[15:0] addr_remain3_247;
address_decode_4 decoder_3_247 = address_decode_4(addr_selector2_15[7],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_247,addr_remain3_247);


wire[15:0] addr_selector3_248;
wire[15:0] addr_remain3_248;
address_decode_4 decoder_3_248 = address_decode_4(addr_selector2_15[8],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_248,addr_remain3_248);


wire[15:0] addr_selector3_249;
wire[15:0] addr_remain3_249;
address_decode_4 decoder_3_249 = address_decode_4(addr_selector2_15[9],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_249,addr_remain3_249);


wire[15:0] addr_selector3_250;
wire[15:0] addr_remain3_250;
address_decode_4 decoder_3_250 = address_decode_4(addr_selector2_15[10],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_250,addr_remain3_250);


wire[15:0] addr_selector3_251;
wire[15:0] addr_remain3_251;
address_decode_4 decoder_3_251 = address_decode_4(addr_selector2_15[11],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_251,addr_remain3_251);


wire[15:0] addr_selector3_252;
wire[15:0] addr_remain3_252;
address_decode_4 decoder_3_252 = address_decode_4(addr_selector2_15[12],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_252,addr_remain3_252);


wire[15:0] addr_selector3_253;
wire[15:0] addr_remain3_253;
address_decode_4 decoder_3_253 = address_decode_4(addr_selector2_15[13],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_253,addr_remain3_253);


wire[15:0] addr_selector3_254;
wire[15:0] addr_remain3_254;
address_decode_4 decoder_3_254 = address_decode_4(addr_selector2_15[14],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_254,addr_remain3_254);


wire[15:0] addr_selector3_255;
wire[15:0] addr_remain3_255;
address_decode_4 decoder_3_255 = address_decode_4(addr_selector2_15[15],addr_remain2_15[15:0],addr_remain2_15,addr_selector3_255,addr_remain3_255);


wire[15:0] addr_selector3_256;
wire[15:0] addr_remain3_256;
address_decode_4 decoder_3_256 = address_decode_4(addr_selector2_16[0],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_256,addr_remain3_256);


wire[15:0] addr_selector3_257;
wire[15:0] addr_remain3_257;
address_decode_4 decoder_3_257 = address_decode_4(addr_selector2_16[1],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_257,addr_remain3_257);


wire[15:0] addr_selector3_258;
wire[15:0] addr_remain3_258;
address_decode_4 decoder_3_258 = address_decode_4(addr_selector2_16[2],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_258,addr_remain3_258);


wire[15:0] addr_selector3_259;
wire[15:0] addr_remain3_259;
address_decode_4 decoder_3_259 = address_decode_4(addr_selector2_16[3],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_259,addr_remain3_259);


wire[15:0] addr_selector3_260;
wire[15:0] addr_remain3_260;
address_decode_4 decoder_3_260 = address_decode_4(addr_selector2_16[4],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_260,addr_remain3_260);


wire[15:0] addr_selector3_261;
wire[15:0] addr_remain3_261;
address_decode_4 decoder_3_261 = address_decode_4(addr_selector2_16[5],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_261,addr_remain3_261);


wire[15:0] addr_selector3_262;
wire[15:0] addr_remain3_262;
address_decode_4 decoder_3_262 = address_decode_4(addr_selector2_16[6],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_262,addr_remain3_262);


wire[15:0] addr_selector3_263;
wire[15:0] addr_remain3_263;
address_decode_4 decoder_3_263 = address_decode_4(addr_selector2_16[7],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_263,addr_remain3_263);


wire[15:0] addr_selector3_264;
wire[15:0] addr_remain3_264;
address_decode_4 decoder_3_264 = address_decode_4(addr_selector2_16[8],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_264,addr_remain3_264);


wire[15:0] addr_selector3_265;
wire[15:0] addr_remain3_265;
address_decode_4 decoder_3_265 = address_decode_4(addr_selector2_16[9],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_265,addr_remain3_265);


wire[15:0] addr_selector3_266;
wire[15:0] addr_remain3_266;
address_decode_4 decoder_3_266 = address_decode_4(addr_selector2_16[10],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_266,addr_remain3_266);


wire[15:0] addr_selector3_267;
wire[15:0] addr_remain3_267;
address_decode_4 decoder_3_267 = address_decode_4(addr_selector2_16[11],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_267,addr_remain3_267);


wire[15:0] addr_selector3_268;
wire[15:0] addr_remain3_268;
address_decode_4 decoder_3_268 = address_decode_4(addr_selector2_16[12],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_268,addr_remain3_268);


wire[15:0] addr_selector3_269;
wire[15:0] addr_remain3_269;
address_decode_4 decoder_3_269 = address_decode_4(addr_selector2_16[13],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_269,addr_remain3_269);


wire[15:0] addr_selector3_270;
wire[15:0] addr_remain3_270;
address_decode_4 decoder_3_270 = address_decode_4(addr_selector2_16[14],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_270,addr_remain3_270);


wire[15:0] addr_selector3_271;
wire[15:0] addr_remain3_271;
address_decode_4 decoder_3_271 = address_decode_4(addr_selector2_16[15],addr_remain2_16[15:0],addr_remain2_16,addr_selector3_271,addr_remain3_271);


wire[15:0] addr_selector3_272;
wire[15:0] addr_remain3_272;
address_decode_4 decoder_3_272 = address_decode_4(addr_selector2_17[0],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_272,addr_remain3_272);


wire[15:0] addr_selector3_273;
wire[15:0] addr_remain3_273;
address_decode_4 decoder_3_273 = address_decode_4(addr_selector2_17[1],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_273,addr_remain3_273);


wire[15:0] addr_selector3_274;
wire[15:0] addr_remain3_274;
address_decode_4 decoder_3_274 = address_decode_4(addr_selector2_17[2],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_274,addr_remain3_274);


wire[15:0] addr_selector3_275;
wire[15:0] addr_remain3_275;
address_decode_4 decoder_3_275 = address_decode_4(addr_selector2_17[3],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_275,addr_remain3_275);


wire[15:0] addr_selector3_276;
wire[15:0] addr_remain3_276;
address_decode_4 decoder_3_276 = address_decode_4(addr_selector2_17[4],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_276,addr_remain3_276);


wire[15:0] addr_selector3_277;
wire[15:0] addr_remain3_277;
address_decode_4 decoder_3_277 = address_decode_4(addr_selector2_17[5],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_277,addr_remain3_277);


wire[15:0] addr_selector3_278;
wire[15:0] addr_remain3_278;
address_decode_4 decoder_3_278 = address_decode_4(addr_selector2_17[6],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_278,addr_remain3_278);


wire[15:0] addr_selector3_279;
wire[15:0] addr_remain3_279;
address_decode_4 decoder_3_279 = address_decode_4(addr_selector2_17[7],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_279,addr_remain3_279);


wire[15:0] addr_selector3_280;
wire[15:0] addr_remain3_280;
address_decode_4 decoder_3_280 = address_decode_4(addr_selector2_17[8],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_280,addr_remain3_280);


wire[15:0] addr_selector3_281;
wire[15:0] addr_remain3_281;
address_decode_4 decoder_3_281 = address_decode_4(addr_selector2_17[9],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_281,addr_remain3_281);


wire[15:0] addr_selector3_282;
wire[15:0] addr_remain3_282;
address_decode_4 decoder_3_282 = address_decode_4(addr_selector2_17[10],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_282,addr_remain3_282);


wire[15:0] addr_selector3_283;
wire[15:0] addr_remain3_283;
address_decode_4 decoder_3_283 = address_decode_4(addr_selector2_17[11],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_283,addr_remain3_283);


wire[15:0] addr_selector3_284;
wire[15:0] addr_remain3_284;
address_decode_4 decoder_3_284 = address_decode_4(addr_selector2_17[12],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_284,addr_remain3_284);


wire[15:0] addr_selector3_285;
wire[15:0] addr_remain3_285;
address_decode_4 decoder_3_285 = address_decode_4(addr_selector2_17[13],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_285,addr_remain3_285);


wire[15:0] addr_selector3_286;
wire[15:0] addr_remain3_286;
address_decode_4 decoder_3_286 = address_decode_4(addr_selector2_17[14],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_286,addr_remain3_286);


wire[15:0] addr_selector3_287;
wire[15:0] addr_remain3_287;
address_decode_4 decoder_3_287 = address_decode_4(addr_selector2_17[15],addr_remain2_17[15:0],addr_remain2_17,addr_selector3_287,addr_remain3_287);


wire[15:0] addr_selector3_288;
wire[15:0] addr_remain3_288;
address_decode_4 decoder_3_288 = address_decode_4(addr_selector2_18[0],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_288,addr_remain3_288);


wire[15:0] addr_selector3_289;
wire[15:0] addr_remain3_289;
address_decode_4 decoder_3_289 = address_decode_4(addr_selector2_18[1],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_289,addr_remain3_289);


wire[15:0] addr_selector3_290;
wire[15:0] addr_remain3_290;
address_decode_4 decoder_3_290 = address_decode_4(addr_selector2_18[2],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_290,addr_remain3_290);


wire[15:0] addr_selector3_291;
wire[15:0] addr_remain3_291;
address_decode_4 decoder_3_291 = address_decode_4(addr_selector2_18[3],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_291,addr_remain3_291);


wire[15:0] addr_selector3_292;
wire[15:0] addr_remain3_292;
address_decode_4 decoder_3_292 = address_decode_4(addr_selector2_18[4],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_292,addr_remain3_292);


wire[15:0] addr_selector3_293;
wire[15:0] addr_remain3_293;
address_decode_4 decoder_3_293 = address_decode_4(addr_selector2_18[5],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_293,addr_remain3_293);


wire[15:0] addr_selector3_294;
wire[15:0] addr_remain3_294;
address_decode_4 decoder_3_294 = address_decode_4(addr_selector2_18[6],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_294,addr_remain3_294);


wire[15:0] addr_selector3_295;
wire[15:0] addr_remain3_295;
address_decode_4 decoder_3_295 = address_decode_4(addr_selector2_18[7],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_295,addr_remain3_295);


wire[15:0] addr_selector3_296;
wire[15:0] addr_remain3_296;
address_decode_4 decoder_3_296 = address_decode_4(addr_selector2_18[8],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_296,addr_remain3_296);


wire[15:0] addr_selector3_297;
wire[15:0] addr_remain3_297;
address_decode_4 decoder_3_297 = address_decode_4(addr_selector2_18[9],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_297,addr_remain3_297);


wire[15:0] addr_selector3_298;
wire[15:0] addr_remain3_298;
address_decode_4 decoder_3_298 = address_decode_4(addr_selector2_18[10],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_298,addr_remain3_298);


wire[15:0] addr_selector3_299;
wire[15:0] addr_remain3_299;
address_decode_4 decoder_3_299 = address_decode_4(addr_selector2_18[11],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_299,addr_remain3_299);


wire[15:0] addr_selector3_300;
wire[15:0] addr_remain3_300;
address_decode_4 decoder_3_300 = address_decode_4(addr_selector2_18[12],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_300,addr_remain3_300);


wire[15:0] addr_selector3_301;
wire[15:0] addr_remain3_301;
address_decode_4 decoder_3_301 = address_decode_4(addr_selector2_18[13],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_301,addr_remain3_301);


wire[15:0] addr_selector3_302;
wire[15:0] addr_remain3_302;
address_decode_4 decoder_3_302 = address_decode_4(addr_selector2_18[14],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_302,addr_remain3_302);


wire[15:0] addr_selector3_303;
wire[15:0] addr_remain3_303;
address_decode_4 decoder_3_303 = address_decode_4(addr_selector2_18[15],addr_remain2_18[15:0],addr_remain2_18,addr_selector3_303,addr_remain3_303);


wire[15:0] addr_selector3_304;
wire[15:0] addr_remain3_304;
address_decode_4 decoder_3_304 = address_decode_4(addr_selector2_19[0],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_304,addr_remain3_304);


wire[15:0] addr_selector3_305;
wire[15:0] addr_remain3_305;
address_decode_4 decoder_3_305 = address_decode_4(addr_selector2_19[1],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_305,addr_remain3_305);


wire[15:0] addr_selector3_306;
wire[15:0] addr_remain3_306;
address_decode_4 decoder_3_306 = address_decode_4(addr_selector2_19[2],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_306,addr_remain3_306);


wire[15:0] addr_selector3_307;
wire[15:0] addr_remain3_307;
address_decode_4 decoder_3_307 = address_decode_4(addr_selector2_19[3],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_307,addr_remain3_307);


wire[15:0] addr_selector3_308;
wire[15:0] addr_remain3_308;
address_decode_4 decoder_3_308 = address_decode_4(addr_selector2_19[4],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_308,addr_remain3_308);


wire[15:0] addr_selector3_309;
wire[15:0] addr_remain3_309;
address_decode_4 decoder_3_309 = address_decode_4(addr_selector2_19[5],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_309,addr_remain3_309);


wire[15:0] addr_selector3_310;
wire[15:0] addr_remain3_310;
address_decode_4 decoder_3_310 = address_decode_4(addr_selector2_19[6],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_310,addr_remain3_310);


wire[15:0] addr_selector3_311;
wire[15:0] addr_remain3_311;
address_decode_4 decoder_3_311 = address_decode_4(addr_selector2_19[7],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_311,addr_remain3_311);


wire[15:0] addr_selector3_312;
wire[15:0] addr_remain3_312;
address_decode_4 decoder_3_312 = address_decode_4(addr_selector2_19[8],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_312,addr_remain3_312);


wire[15:0] addr_selector3_313;
wire[15:0] addr_remain3_313;
address_decode_4 decoder_3_313 = address_decode_4(addr_selector2_19[9],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_313,addr_remain3_313);


wire[15:0] addr_selector3_314;
wire[15:0] addr_remain3_314;
address_decode_4 decoder_3_314 = address_decode_4(addr_selector2_19[10],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_314,addr_remain3_314);


wire[15:0] addr_selector3_315;
wire[15:0] addr_remain3_315;
address_decode_4 decoder_3_315 = address_decode_4(addr_selector2_19[11],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_315,addr_remain3_315);


wire[15:0] addr_selector3_316;
wire[15:0] addr_remain3_316;
address_decode_4 decoder_3_316 = address_decode_4(addr_selector2_19[12],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_316,addr_remain3_316);


wire[15:0] addr_selector3_317;
wire[15:0] addr_remain3_317;
address_decode_4 decoder_3_317 = address_decode_4(addr_selector2_19[13],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_317,addr_remain3_317);


wire[15:0] addr_selector3_318;
wire[15:0] addr_remain3_318;
address_decode_4 decoder_3_318 = address_decode_4(addr_selector2_19[14],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_318,addr_remain3_318);


wire[15:0] addr_selector3_319;
wire[15:0] addr_remain3_319;
address_decode_4 decoder_3_319 = address_decode_4(addr_selector2_19[15],addr_remain2_19[15:0],addr_remain2_19,addr_selector3_319,addr_remain3_319);


wire[15:0] addr_selector3_320;
wire[15:0] addr_remain3_320;
address_decode_4 decoder_3_320 = address_decode_4(addr_selector2_20[0],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_320,addr_remain3_320);


wire[15:0] addr_selector3_321;
wire[15:0] addr_remain3_321;
address_decode_4 decoder_3_321 = address_decode_4(addr_selector2_20[1],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_321,addr_remain3_321);


wire[15:0] addr_selector3_322;
wire[15:0] addr_remain3_322;
address_decode_4 decoder_3_322 = address_decode_4(addr_selector2_20[2],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_322,addr_remain3_322);


wire[15:0] addr_selector3_323;
wire[15:0] addr_remain3_323;
address_decode_4 decoder_3_323 = address_decode_4(addr_selector2_20[3],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_323,addr_remain3_323);


wire[15:0] addr_selector3_324;
wire[15:0] addr_remain3_324;
address_decode_4 decoder_3_324 = address_decode_4(addr_selector2_20[4],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_324,addr_remain3_324);


wire[15:0] addr_selector3_325;
wire[15:0] addr_remain3_325;
address_decode_4 decoder_3_325 = address_decode_4(addr_selector2_20[5],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_325,addr_remain3_325);


wire[15:0] addr_selector3_326;
wire[15:0] addr_remain3_326;
address_decode_4 decoder_3_326 = address_decode_4(addr_selector2_20[6],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_326,addr_remain3_326);


wire[15:0] addr_selector3_327;
wire[15:0] addr_remain3_327;
address_decode_4 decoder_3_327 = address_decode_4(addr_selector2_20[7],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_327,addr_remain3_327);


wire[15:0] addr_selector3_328;
wire[15:0] addr_remain3_328;
address_decode_4 decoder_3_328 = address_decode_4(addr_selector2_20[8],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_328,addr_remain3_328);


wire[15:0] addr_selector3_329;
wire[15:0] addr_remain3_329;
address_decode_4 decoder_3_329 = address_decode_4(addr_selector2_20[9],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_329,addr_remain3_329);


wire[15:0] addr_selector3_330;
wire[15:0] addr_remain3_330;
address_decode_4 decoder_3_330 = address_decode_4(addr_selector2_20[10],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_330,addr_remain3_330);


wire[15:0] addr_selector3_331;
wire[15:0] addr_remain3_331;
address_decode_4 decoder_3_331 = address_decode_4(addr_selector2_20[11],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_331,addr_remain3_331);


wire[15:0] addr_selector3_332;
wire[15:0] addr_remain3_332;
address_decode_4 decoder_3_332 = address_decode_4(addr_selector2_20[12],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_332,addr_remain3_332);


wire[15:0] addr_selector3_333;
wire[15:0] addr_remain3_333;
address_decode_4 decoder_3_333 = address_decode_4(addr_selector2_20[13],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_333,addr_remain3_333);


wire[15:0] addr_selector3_334;
wire[15:0] addr_remain3_334;
address_decode_4 decoder_3_334 = address_decode_4(addr_selector2_20[14],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_334,addr_remain3_334);


wire[15:0] addr_selector3_335;
wire[15:0] addr_remain3_335;
address_decode_4 decoder_3_335 = address_decode_4(addr_selector2_20[15],addr_remain2_20[15:0],addr_remain2_20,addr_selector3_335,addr_remain3_335);


wire[15:0] addr_selector3_336;
wire[15:0] addr_remain3_336;
address_decode_4 decoder_3_336 = address_decode_4(addr_selector2_21[0],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_336,addr_remain3_336);


wire[15:0] addr_selector3_337;
wire[15:0] addr_remain3_337;
address_decode_4 decoder_3_337 = address_decode_4(addr_selector2_21[1],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_337,addr_remain3_337);


wire[15:0] addr_selector3_338;
wire[15:0] addr_remain3_338;
address_decode_4 decoder_3_338 = address_decode_4(addr_selector2_21[2],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_338,addr_remain3_338);


wire[15:0] addr_selector3_339;
wire[15:0] addr_remain3_339;
address_decode_4 decoder_3_339 = address_decode_4(addr_selector2_21[3],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_339,addr_remain3_339);


wire[15:0] addr_selector3_340;
wire[15:0] addr_remain3_340;
address_decode_4 decoder_3_340 = address_decode_4(addr_selector2_21[4],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_340,addr_remain3_340);


wire[15:0] addr_selector3_341;
wire[15:0] addr_remain3_341;
address_decode_4 decoder_3_341 = address_decode_4(addr_selector2_21[5],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_341,addr_remain3_341);


wire[15:0] addr_selector3_342;
wire[15:0] addr_remain3_342;
address_decode_4 decoder_3_342 = address_decode_4(addr_selector2_21[6],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_342,addr_remain3_342);


wire[15:0] addr_selector3_343;
wire[15:0] addr_remain3_343;
address_decode_4 decoder_3_343 = address_decode_4(addr_selector2_21[7],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_343,addr_remain3_343);


wire[15:0] addr_selector3_344;
wire[15:0] addr_remain3_344;
address_decode_4 decoder_3_344 = address_decode_4(addr_selector2_21[8],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_344,addr_remain3_344);


wire[15:0] addr_selector3_345;
wire[15:0] addr_remain3_345;
address_decode_4 decoder_3_345 = address_decode_4(addr_selector2_21[9],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_345,addr_remain3_345);


wire[15:0] addr_selector3_346;
wire[15:0] addr_remain3_346;
address_decode_4 decoder_3_346 = address_decode_4(addr_selector2_21[10],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_346,addr_remain3_346);


wire[15:0] addr_selector3_347;
wire[15:0] addr_remain3_347;
address_decode_4 decoder_3_347 = address_decode_4(addr_selector2_21[11],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_347,addr_remain3_347);


wire[15:0] addr_selector3_348;
wire[15:0] addr_remain3_348;
address_decode_4 decoder_3_348 = address_decode_4(addr_selector2_21[12],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_348,addr_remain3_348);


wire[15:0] addr_selector3_349;
wire[15:0] addr_remain3_349;
address_decode_4 decoder_3_349 = address_decode_4(addr_selector2_21[13],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_349,addr_remain3_349);


wire[15:0] addr_selector3_350;
wire[15:0] addr_remain3_350;
address_decode_4 decoder_3_350 = address_decode_4(addr_selector2_21[14],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_350,addr_remain3_350);


wire[15:0] addr_selector3_351;
wire[15:0] addr_remain3_351;
address_decode_4 decoder_3_351 = address_decode_4(addr_selector2_21[15],addr_remain2_21[15:0],addr_remain2_21,addr_selector3_351,addr_remain3_351);


wire[15:0] addr_selector3_352;
wire[15:0] addr_remain3_352;
address_decode_4 decoder_3_352 = address_decode_4(addr_selector2_22[0],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_352,addr_remain3_352);


wire[15:0] addr_selector3_353;
wire[15:0] addr_remain3_353;
address_decode_4 decoder_3_353 = address_decode_4(addr_selector2_22[1],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_353,addr_remain3_353);


wire[15:0] addr_selector3_354;
wire[15:0] addr_remain3_354;
address_decode_4 decoder_3_354 = address_decode_4(addr_selector2_22[2],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_354,addr_remain3_354);


wire[15:0] addr_selector3_355;
wire[15:0] addr_remain3_355;
address_decode_4 decoder_3_355 = address_decode_4(addr_selector2_22[3],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_355,addr_remain3_355);


wire[15:0] addr_selector3_356;
wire[15:0] addr_remain3_356;
address_decode_4 decoder_3_356 = address_decode_4(addr_selector2_22[4],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_356,addr_remain3_356);


wire[15:0] addr_selector3_357;
wire[15:0] addr_remain3_357;
address_decode_4 decoder_3_357 = address_decode_4(addr_selector2_22[5],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_357,addr_remain3_357);


wire[15:0] addr_selector3_358;
wire[15:0] addr_remain3_358;
address_decode_4 decoder_3_358 = address_decode_4(addr_selector2_22[6],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_358,addr_remain3_358);


wire[15:0] addr_selector3_359;
wire[15:0] addr_remain3_359;
address_decode_4 decoder_3_359 = address_decode_4(addr_selector2_22[7],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_359,addr_remain3_359);


wire[15:0] addr_selector3_360;
wire[15:0] addr_remain3_360;
address_decode_4 decoder_3_360 = address_decode_4(addr_selector2_22[8],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_360,addr_remain3_360);


wire[15:0] addr_selector3_361;
wire[15:0] addr_remain3_361;
address_decode_4 decoder_3_361 = address_decode_4(addr_selector2_22[9],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_361,addr_remain3_361);


wire[15:0] addr_selector3_362;
wire[15:0] addr_remain3_362;
address_decode_4 decoder_3_362 = address_decode_4(addr_selector2_22[10],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_362,addr_remain3_362);


wire[15:0] addr_selector3_363;
wire[15:0] addr_remain3_363;
address_decode_4 decoder_3_363 = address_decode_4(addr_selector2_22[11],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_363,addr_remain3_363);


wire[15:0] addr_selector3_364;
wire[15:0] addr_remain3_364;
address_decode_4 decoder_3_364 = address_decode_4(addr_selector2_22[12],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_364,addr_remain3_364);


wire[15:0] addr_selector3_365;
wire[15:0] addr_remain3_365;
address_decode_4 decoder_3_365 = address_decode_4(addr_selector2_22[13],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_365,addr_remain3_365);


wire[15:0] addr_selector3_366;
wire[15:0] addr_remain3_366;
address_decode_4 decoder_3_366 = address_decode_4(addr_selector2_22[14],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_366,addr_remain3_366);


wire[15:0] addr_selector3_367;
wire[15:0] addr_remain3_367;
address_decode_4 decoder_3_367 = address_decode_4(addr_selector2_22[15],addr_remain2_22[15:0],addr_remain2_22,addr_selector3_367,addr_remain3_367);


wire[15:0] addr_selector3_368;
wire[15:0] addr_remain3_368;
address_decode_4 decoder_3_368 = address_decode_4(addr_selector2_23[0],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_368,addr_remain3_368);


wire[15:0] addr_selector3_369;
wire[15:0] addr_remain3_369;
address_decode_4 decoder_3_369 = address_decode_4(addr_selector2_23[1],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_369,addr_remain3_369);


wire[15:0] addr_selector3_370;
wire[15:0] addr_remain3_370;
address_decode_4 decoder_3_370 = address_decode_4(addr_selector2_23[2],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_370,addr_remain3_370);


wire[15:0] addr_selector3_371;
wire[15:0] addr_remain3_371;
address_decode_4 decoder_3_371 = address_decode_4(addr_selector2_23[3],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_371,addr_remain3_371);


wire[15:0] addr_selector3_372;
wire[15:0] addr_remain3_372;
address_decode_4 decoder_3_372 = address_decode_4(addr_selector2_23[4],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_372,addr_remain3_372);


wire[15:0] addr_selector3_373;
wire[15:0] addr_remain3_373;
address_decode_4 decoder_3_373 = address_decode_4(addr_selector2_23[5],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_373,addr_remain3_373);


wire[15:0] addr_selector3_374;
wire[15:0] addr_remain3_374;
address_decode_4 decoder_3_374 = address_decode_4(addr_selector2_23[6],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_374,addr_remain3_374);


wire[15:0] addr_selector3_375;
wire[15:0] addr_remain3_375;
address_decode_4 decoder_3_375 = address_decode_4(addr_selector2_23[7],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_375,addr_remain3_375);


wire[15:0] addr_selector3_376;
wire[15:0] addr_remain3_376;
address_decode_4 decoder_3_376 = address_decode_4(addr_selector2_23[8],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_376,addr_remain3_376);


wire[15:0] addr_selector3_377;
wire[15:0] addr_remain3_377;
address_decode_4 decoder_3_377 = address_decode_4(addr_selector2_23[9],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_377,addr_remain3_377);


wire[15:0] addr_selector3_378;
wire[15:0] addr_remain3_378;
address_decode_4 decoder_3_378 = address_decode_4(addr_selector2_23[10],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_378,addr_remain3_378);


wire[15:0] addr_selector3_379;
wire[15:0] addr_remain3_379;
address_decode_4 decoder_3_379 = address_decode_4(addr_selector2_23[11],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_379,addr_remain3_379);


wire[15:0] addr_selector3_380;
wire[15:0] addr_remain3_380;
address_decode_4 decoder_3_380 = address_decode_4(addr_selector2_23[12],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_380,addr_remain3_380);


wire[15:0] addr_selector3_381;
wire[15:0] addr_remain3_381;
address_decode_4 decoder_3_381 = address_decode_4(addr_selector2_23[13],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_381,addr_remain3_381);


wire[15:0] addr_selector3_382;
wire[15:0] addr_remain3_382;
address_decode_4 decoder_3_382 = address_decode_4(addr_selector2_23[14],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_382,addr_remain3_382);


wire[15:0] addr_selector3_383;
wire[15:0] addr_remain3_383;
address_decode_4 decoder_3_383 = address_decode_4(addr_selector2_23[15],addr_remain2_23[15:0],addr_remain2_23,addr_selector3_383,addr_remain3_383);


wire[15:0] addr_selector3_384;
wire[15:0] addr_remain3_384;
address_decode_4 decoder_3_384 = address_decode_4(addr_selector2_24[0],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_384,addr_remain3_384);


wire[15:0] addr_selector3_385;
wire[15:0] addr_remain3_385;
address_decode_4 decoder_3_385 = address_decode_4(addr_selector2_24[1],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_385,addr_remain3_385);


wire[15:0] addr_selector3_386;
wire[15:0] addr_remain3_386;
address_decode_4 decoder_3_386 = address_decode_4(addr_selector2_24[2],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_386,addr_remain3_386);


wire[15:0] addr_selector3_387;
wire[15:0] addr_remain3_387;
address_decode_4 decoder_3_387 = address_decode_4(addr_selector2_24[3],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_387,addr_remain3_387);


wire[15:0] addr_selector3_388;
wire[15:0] addr_remain3_388;
address_decode_4 decoder_3_388 = address_decode_4(addr_selector2_24[4],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_388,addr_remain3_388);


wire[15:0] addr_selector3_389;
wire[15:0] addr_remain3_389;
address_decode_4 decoder_3_389 = address_decode_4(addr_selector2_24[5],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_389,addr_remain3_389);


wire[15:0] addr_selector3_390;
wire[15:0] addr_remain3_390;
address_decode_4 decoder_3_390 = address_decode_4(addr_selector2_24[6],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_390,addr_remain3_390);


wire[15:0] addr_selector3_391;
wire[15:0] addr_remain3_391;
address_decode_4 decoder_3_391 = address_decode_4(addr_selector2_24[7],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_391,addr_remain3_391);


wire[15:0] addr_selector3_392;
wire[15:0] addr_remain3_392;
address_decode_4 decoder_3_392 = address_decode_4(addr_selector2_24[8],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_392,addr_remain3_392);


wire[15:0] addr_selector3_393;
wire[15:0] addr_remain3_393;
address_decode_4 decoder_3_393 = address_decode_4(addr_selector2_24[9],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_393,addr_remain3_393);


wire[15:0] addr_selector3_394;
wire[15:0] addr_remain3_394;
address_decode_4 decoder_3_394 = address_decode_4(addr_selector2_24[10],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_394,addr_remain3_394);


wire[15:0] addr_selector3_395;
wire[15:0] addr_remain3_395;
address_decode_4 decoder_3_395 = address_decode_4(addr_selector2_24[11],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_395,addr_remain3_395);


wire[15:0] addr_selector3_396;
wire[15:0] addr_remain3_396;
address_decode_4 decoder_3_396 = address_decode_4(addr_selector2_24[12],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_396,addr_remain3_396);


wire[15:0] addr_selector3_397;
wire[15:0] addr_remain3_397;
address_decode_4 decoder_3_397 = address_decode_4(addr_selector2_24[13],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_397,addr_remain3_397);


wire[15:0] addr_selector3_398;
wire[15:0] addr_remain3_398;
address_decode_4 decoder_3_398 = address_decode_4(addr_selector2_24[14],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_398,addr_remain3_398);


wire[15:0] addr_selector3_399;
wire[15:0] addr_remain3_399;
address_decode_4 decoder_3_399 = address_decode_4(addr_selector2_24[15],addr_remain2_24[15:0],addr_remain2_24,addr_selector3_399,addr_remain3_399);


wire[15:0] addr_selector3_400;
wire[15:0] addr_remain3_400;
address_decode_4 decoder_3_400 = address_decode_4(addr_selector2_25[0],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_400,addr_remain3_400);


wire[15:0] addr_selector3_401;
wire[15:0] addr_remain3_401;
address_decode_4 decoder_3_401 = address_decode_4(addr_selector2_25[1],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_401,addr_remain3_401);


wire[15:0] addr_selector3_402;
wire[15:0] addr_remain3_402;
address_decode_4 decoder_3_402 = address_decode_4(addr_selector2_25[2],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_402,addr_remain3_402);


wire[15:0] addr_selector3_403;
wire[15:0] addr_remain3_403;
address_decode_4 decoder_3_403 = address_decode_4(addr_selector2_25[3],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_403,addr_remain3_403);


wire[15:0] addr_selector3_404;
wire[15:0] addr_remain3_404;
address_decode_4 decoder_3_404 = address_decode_4(addr_selector2_25[4],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_404,addr_remain3_404);


wire[15:0] addr_selector3_405;
wire[15:0] addr_remain3_405;
address_decode_4 decoder_3_405 = address_decode_4(addr_selector2_25[5],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_405,addr_remain3_405);


wire[15:0] addr_selector3_406;
wire[15:0] addr_remain3_406;
address_decode_4 decoder_3_406 = address_decode_4(addr_selector2_25[6],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_406,addr_remain3_406);


wire[15:0] addr_selector3_407;
wire[15:0] addr_remain3_407;
address_decode_4 decoder_3_407 = address_decode_4(addr_selector2_25[7],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_407,addr_remain3_407);


wire[15:0] addr_selector3_408;
wire[15:0] addr_remain3_408;
address_decode_4 decoder_3_408 = address_decode_4(addr_selector2_25[8],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_408,addr_remain3_408);


wire[15:0] addr_selector3_409;
wire[15:0] addr_remain3_409;
address_decode_4 decoder_3_409 = address_decode_4(addr_selector2_25[9],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_409,addr_remain3_409);


wire[15:0] addr_selector3_410;
wire[15:0] addr_remain3_410;
address_decode_4 decoder_3_410 = address_decode_4(addr_selector2_25[10],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_410,addr_remain3_410);


wire[15:0] addr_selector3_411;
wire[15:0] addr_remain3_411;
address_decode_4 decoder_3_411 = address_decode_4(addr_selector2_25[11],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_411,addr_remain3_411);


wire[15:0] addr_selector3_412;
wire[15:0] addr_remain3_412;
address_decode_4 decoder_3_412 = address_decode_4(addr_selector2_25[12],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_412,addr_remain3_412);


wire[15:0] addr_selector3_413;
wire[15:0] addr_remain3_413;
address_decode_4 decoder_3_413 = address_decode_4(addr_selector2_25[13],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_413,addr_remain3_413);


wire[15:0] addr_selector3_414;
wire[15:0] addr_remain3_414;
address_decode_4 decoder_3_414 = address_decode_4(addr_selector2_25[14],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_414,addr_remain3_414);


wire[15:0] addr_selector3_415;
wire[15:0] addr_remain3_415;
address_decode_4 decoder_3_415 = address_decode_4(addr_selector2_25[15],addr_remain2_25[15:0],addr_remain2_25,addr_selector3_415,addr_remain3_415);


wire[15:0] addr_selector3_416;
wire[15:0] addr_remain3_416;
address_decode_4 decoder_3_416 = address_decode_4(addr_selector2_26[0],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_416,addr_remain3_416);


wire[15:0] addr_selector3_417;
wire[15:0] addr_remain3_417;
address_decode_4 decoder_3_417 = address_decode_4(addr_selector2_26[1],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_417,addr_remain3_417);


wire[15:0] addr_selector3_418;
wire[15:0] addr_remain3_418;
address_decode_4 decoder_3_418 = address_decode_4(addr_selector2_26[2],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_418,addr_remain3_418);


wire[15:0] addr_selector3_419;
wire[15:0] addr_remain3_419;
address_decode_4 decoder_3_419 = address_decode_4(addr_selector2_26[3],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_419,addr_remain3_419);


wire[15:0] addr_selector3_420;
wire[15:0] addr_remain3_420;
address_decode_4 decoder_3_420 = address_decode_4(addr_selector2_26[4],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_420,addr_remain3_420);


wire[15:0] addr_selector3_421;
wire[15:0] addr_remain3_421;
address_decode_4 decoder_3_421 = address_decode_4(addr_selector2_26[5],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_421,addr_remain3_421);


wire[15:0] addr_selector3_422;
wire[15:0] addr_remain3_422;
address_decode_4 decoder_3_422 = address_decode_4(addr_selector2_26[6],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_422,addr_remain3_422);


wire[15:0] addr_selector3_423;
wire[15:0] addr_remain3_423;
address_decode_4 decoder_3_423 = address_decode_4(addr_selector2_26[7],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_423,addr_remain3_423);


wire[15:0] addr_selector3_424;
wire[15:0] addr_remain3_424;
address_decode_4 decoder_3_424 = address_decode_4(addr_selector2_26[8],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_424,addr_remain3_424);


wire[15:0] addr_selector3_425;
wire[15:0] addr_remain3_425;
address_decode_4 decoder_3_425 = address_decode_4(addr_selector2_26[9],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_425,addr_remain3_425);


wire[15:0] addr_selector3_426;
wire[15:0] addr_remain3_426;
address_decode_4 decoder_3_426 = address_decode_4(addr_selector2_26[10],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_426,addr_remain3_426);


wire[15:0] addr_selector3_427;
wire[15:0] addr_remain3_427;
address_decode_4 decoder_3_427 = address_decode_4(addr_selector2_26[11],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_427,addr_remain3_427);


wire[15:0] addr_selector3_428;
wire[15:0] addr_remain3_428;
address_decode_4 decoder_3_428 = address_decode_4(addr_selector2_26[12],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_428,addr_remain3_428);


wire[15:0] addr_selector3_429;
wire[15:0] addr_remain3_429;
address_decode_4 decoder_3_429 = address_decode_4(addr_selector2_26[13],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_429,addr_remain3_429);


wire[15:0] addr_selector3_430;
wire[15:0] addr_remain3_430;
address_decode_4 decoder_3_430 = address_decode_4(addr_selector2_26[14],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_430,addr_remain3_430);


wire[15:0] addr_selector3_431;
wire[15:0] addr_remain3_431;
address_decode_4 decoder_3_431 = address_decode_4(addr_selector2_26[15],addr_remain2_26[15:0],addr_remain2_26,addr_selector3_431,addr_remain3_431);


wire[15:0] addr_selector3_432;
wire[15:0] addr_remain3_432;
address_decode_4 decoder_3_432 = address_decode_4(addr_selector2_27[0],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_432,addr_remain3_432);


wire[15:0] addr_selector3_433;
wire[15:0] addr_remain3_433;
address_decode_4 decoder_3_433 = address_decode_4(addr_selector2_27[1],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_433,addr_remain3_433);


wire[15:0] addr_selector3_434;
wire[15:0] addr_remain3_434;
address_decode_4 decoder_3_434 = address_decode_4(addr_selector2_27[2],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_434,addr_remain3_434);


wire[15:0] addr_selector3_435;
wire[15:0] addr_remain3_435;
address_decode_4 decoder_3_435 = address_decode_4(addr_selector2_27[3],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_435,addr_remain3_435);


wire[15:0] addr_selector3_436;
wire[15:0] addr_remain3_436;
address_decode_4 decoder_3_436 = address_decode_4(addr_selector2_27[4],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_436,addr_remain3_436);


wire[15:0] addr_selector3_437;
wire[15:0] addr_remain3_437;
address_decode_4 decoder_3_437 = address_decode_4(addr_selector2_27[5],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_437,addr_remain3_437);


wire[15:0] addr_selector3_438;
wire[15:0] addr_remain3_438;
address_decode_4 decoder_3_438 = address_decode_4(addr_selector2_27[6],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_438,addr_remain3_438);


wire[15:0] addr_selector3_439;
wire[15:0] addr_remain3_439;
address_decode_4 decoder_3_439 = address_decode_4(addr_selector2_27[7],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_439,addr_remain3_439);


wire[15:0] addr_selector3_440;
wire[15:0] addr_remain3_440;
address_decode_4 decoder_3_440 = address_decode_4(addr_selector2_27[8],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_440,addr_remain3_440);


wire[15:0] addr_selector3_441;
wire[15:0] addr_remain3_441;
address_decode_4 decoder_3_441 = address_decode_4(addr_selector2_27[9],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_441,addr_remain3_441);


wire[15:0] addr_selector3_442;
wire[15:0] addr_remain3_442;
address_decode_4 decoder_3_442 = address_decode_4(addr_selector2_27[10],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_442,addr_remain3_442);


wire[15:0] addr_selector3_443;
wire[15:0] addr_remain3_443;
address_decode_4 decoder_3_443 = address_decode_4(addr_selector2_27[11],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_443,addr_remain3_443);


wire[15:0] addr_selector3_444;
wire[15:0] addr_remain3_444;
address_decode_4 decoder_3_444 = address_decode_4(addr_selector2_27[12],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_444,addr_remain3_444);


wire[15:0] addr_selector3_445;
wire[15:0] addr_remain3_445;
address_decode_4 decoder_3_445 = address_decode_4(addr_selector2_27[13],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_445,addr_remain3_445);


wire[15:0] addr_selector3_446;
wire[15:0] addr_remain3_446;
address_decode_4 decoder_3_446 = address_decode_4(addr_selector2_27[14],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_446,addr_remain3_446);


wire[15:0] addr_selector3_447;
wire[15:0] addr_remain3_447;
address_decode_4 decoder_3_447 = address_decode_4(addr_selector2_27[15],addr_remain2_27[15:0],addr_remain2_27,addr_selector3_447,addr_remain3_447);


wire[15:0] addr_selector3_448;
wire[15:0] addr_remain3_448;
address_decode_4 decoder_3_448 = address_decode_4(addr_selector2_28[0],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_448,addr_remain3_448);


wire[15:0] addr_selector3_449;
wire[15:0] addr_remain3_449;
address_decode_4 decoder_3_449 = address_decode_4(addr_selector2_28[1],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_449,addr_remain3_449);


wire[15:0] addr_selector3_450;
wire[15:0] addr_remain3_450;
address_decode_4 decoder_3_450 = address_decode_4(addr_selector2_28[2],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_450,addr_remain3_450);


wire[15:0] addr_selector3_451;
wire[15:0] addr_remain3_451;
address_decode_4 decoder_3_451 = address_decode_4(addr_selector2_28[3],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_451,addr_remain3_451);


wire[15:0] addr_selector3_452;
wire[15:0] addr_remain3_452;
address_decode_4 decoder_3_452 = address_decode_4(addr_selector2_28[4],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_452,addr_remain3_452);


wire[15:0] addr_selector3_453;
wire[15:0] addr_remain3_453;
address_decode_4 decoder_3_453 = address_decode_4(addr_selector2_28[5],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_453,addr_remain3_453);


wire[15:0] addr_selector3_454;
wire[15:0] addr_remain3_454;
address_decode_4 decoder_3_454 = address_decode_4(addr_selector2_28[6],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_454,addr_remain3_454);


wire[15:0] addr_selector3_455;
wire[15:0] addr_remain3_455;
address_decode_4 decoder_3_455 = address_decode_4(addr_selector2_28[7],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_455,addr_remain3_455);


wire[15:0] addr_selector3_456;
wire[15:0] addr_remain3_456;
address_decode_4 decoder_3_456 = address_decode_4(addr_selector2_28[8],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_456,addr_remain3_456);


wire[15:0] addr_selector3_457;
wire[15:0] addr_remain3_457;
address_decode_4 decoder_3_457 = address_decode_4(addr_selector2_28[9],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_457,addr_remain3_457);


wire[15:0] addr_selector3_458;
wire[15:0] addr_remain3_458;
address_decode_4 decoder_3_458 = address_decode_4(addr_selector2_28[10],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_458,addr_remain3_458);


wire[15:0] addr_selector3_459;
wire[15:0] addr_remain3_459;
address_decode_4 decoder_3_459 = address_decode_4(addr_selector2_28[11],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_459,addr_remain3_459);


wire[15:0] addr_selector3_460;
wire[15:0] addr_remain3_460;
address_decode_4 decoder_3_460 = address_decode_4(addr_selector2_28[12],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_460,addr_remain3_460);


wire[15:0] addr_selector3_461;
wire[15:0] addr_remain3_461;
address_decode_4 decoder_3_461 = address_decode_4(addr_selector2_28[13],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_461,addr_remain3_461);


wire[15:0] addr_selector3_462;
wire[15:0] addr_remain3_462;
address_decode_4 decoder_3_462 = address_decode_4(addr_selector2_28[14],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_462,addr_remain3_462);


wire[15:0] addr_selector3_463;
wire[15:0] addr_remain3_463;
address_decode_4 decoder_3_463 = address_decode_4(addr_selector2_28[15],addr_remain2_28[15:0],addr_remain2_28,addr_selector3_463,addr_remain3_463);


wire[15:0] addr_selector3_464;
wire[15:0] addr_remain3_464;
address_decode_4 decoder_3_464 = address_decode_4(addr_selector2_29[0],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_464,addr_remain3_464);


wire[15:0] addr_selector3_465;
wire[15:0] addr_remain3_465;
address_decode_4 decoder_3_465 = address_decode_4(addr_selector2_29[1],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_465,addr_remain3_465);


wire[15:0] addr_selector3_466;
wire[15:0] addr_remain3_466;
address_decode_4 decoder_3_466 = address_decode_4(addr_selector2_29[2],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_466,addr_remain3_466);


wire[15:0] addr_selector3_467;
wire[15:0] addr_remain3_467;
address_decode_4 decoder_3_467 = address_decode_4(addr_selector2_29[3],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_467,addr_remain3_467);


wire[15:0] addr_selector3_468;
wire[15:0] addr_remain3_468;
address_decode_4 decoder_3_468 = address_decode_4(addr_selector2_29[4],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_468,addr_remain3_468);


wire[15:0] addr_selector3_469;
wire[15:0] addr_remain3_469;
address_decode_4 decoder_3_469 = address_decode_4(addr_selector2_29[5],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_469,addr_remain3_469);


wire[15:0] addr_selector3_470;
wire[15:0] addr_remain3_470;
address_decode_4 decoder_3_470 = address_decode_4(addr_selector2_29[6],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_470,addr_remain3_470);


wire[15:0] addr_selector3_471;
wire[15:0] addr_remain3_471;
address_decode_4 decoder_3_471 = address_decode_4(addr_selector2_29[7],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_471,addr_remain3_471);


wire[15:0] addr_selector3_472;
wire[15:0] addr_remain3_472;
address_decode_4 decoder_3_472 = address_decode_4(addr_selector2_29[8],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_472,addr_remain3_472);


wire[15:0] addr_selector3_473;
wire[15:0] addr_remain3_473;
address_decode_4 decoder_3_473 = address_decode_4(addr_selector2_29[9],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_473,addr_remain3_473);


wire[15:0] addr_selector3_474;
wire[15:0] addr_remain3_474;
address_decode_4 decoder_3_474 = address_decode_4(addr_selector2_29[10],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_474,addr_remain3_474);


wire[15:0] addr_selector3_475;
wire[15:0] addr_remain3_475;
address_decode_4 decoder_3_475 = address_decode_4(addr_selector2_29[11],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_475,addr_remain3_475);


wire[15:0] addr_selector3_476;
wire[15:0] addr_remain3_476;
address_decode_4 decoder_3_476 = address_decode_4(addr_selector2_29[12],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_476,addr_remain3_476);


wire[15:0] addr_selector3_477;
wire[15:0] addr_remain3_477;
address_decode_4 decoder_3_477 = address_decode_4(addr_selector2_29[13],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_477,addr_remain3_477);


wire[15:0] addr_selector3_478;
wire[15:0] addr_remain3_478;
address_decode_4 decoder_3_478 = address_decode_4(addr_selector2_29[14],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_478,addr_remain3_478);


wire[15:0] addr_selector3_479;
wire[15:0] addr_remain3_479;
address_decode_4 decoder_3_479 = address_decode_4(addr_selector2_29[15],addr_remain2_29[15:0],addr_remain2_29,addr_selector3_479,addr_remain3_479);


wire[15:0] addr_selector3_480;
wire[15:0] addr_remain3_480;
address_decode_4 decoder_3_480 = address_decode_4(addr_selector2_30[0],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_480,addr_remain3_480);


wire[15:0] addr_selector3_481;
wire[15:0] addr_remain3_481;
address_decode_4 decoder_3_481 = address_decode_4(addr_selector2_30[1],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_481,addr_remain3_481);


wire[15:0] addr_selector3_482;
wire[15:0] addr_remain3_482;
address_decode_4 decoder_3_482 = address_decode_4(addr_selector2_30[2],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_482,addr_remain3_482);


wire[15:0] addr_selector3_483;
wire[15:0] addr_remain3_483;
address_decode_4 decoder_3_483 = address_decode_4(addr_selector2_30[3],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_483,addr_remain3_483);


wire[15:0] addr_selector3_484;
wire[15:0] addr_remain3_484;
address_decode_4 decoder_3_484 = address_decode_4(addr_selector2_30[4],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_484,addr_remain3_484);


wire[15:0] addr_selector3_485;
wire[15:0] addr_remain3_485;
address_decode_4 decoder_3_485 = address_decode_4(addr_selector2_30[5],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_485,addr_remain3_485);


wire[15:0] addr_selector3_486;
wire[15:0] addr_remain3_486;
address_decode_4 decoder_3_486 = address_decode_4(addr_selector2_30[6],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_486,addr_remain3_486);


wire[15:0] addr_selector3_487;
wire[15:0] addr_remain3_487;
address_decode_4 decoder_3_487 = address_decode_4(addr_selector2_30[7],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_487,addr_remain3_487);


wire[15:0] addr_selector3_488;
wire[15:0] addr_remain3_488;
address_decode_4 decoder_3_488 = address_decode_4(addr_selector2_30[8],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_488,addr_remain3_488);


wire[15:0] addr_selector3_489;
wire[15:0] addr_remain3_489;
address_decode_4 decoder_3_489 = address_decode_4(addr_selector2_30[9],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_489,addr_remain3_489);


wire[15:0] addr_selector3_490;
wire[15:0] addr_remain3_490;
address_decode_4 decoder_3_490 = address_decode_4(addr_selector2_30[10],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_490,addr_remain3_490);


wire[15:0] addr_selector3_491;
wire[15:0] addr_remain3_491;
address_decode_4 decoder_3_491 = address_decode_4(addr_selector2_30[11],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_491,addr_remain3_491);


wire[15:0] addr_selector3_492;
wire[15:0] addr_remain3_492;
address_decode_4 decoder_3_492 = address_decode_4(addr_selector2_30[12],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_492,addr_remain3_492);


wire[15:0] addr_selector3_493;
wire[15:0] addr_remain3_493;
address_decode_4 decoder_3_493 = address_decode_4(addr_selector2_30[13],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_493,addr_remain3_493);


wire[15:0] addr_selector3_494;
wire[15:0] addr_remain3_494;
address_decode_4 decoder_3_494 = address_decode_4(addr_selector2_30[14],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_494,addr_remain3_494);


wire[15:0] addr_selector3_495;
wire[15:0] addr_remain3_495;
address_decode_4 decoder_3_495 = address_decode_4(addr_selector2_30[15],addr_remain2_30[15:0],addr_remain2_30,addr_selector3_495,addr_remain3_495);


wire[15:0] addr_selector3_496;
wire[15:0] addr_remain3_496;
address_decode_4 decoder_3_496 = address_decode_4(addr_selector2_31[0],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_496,addr_remain3_496);


wire[15:0] addr_selector3_497;
wire[15:0] addr_remain3_497;
address_decode_4 decoder_3_497 = address_decode_4(addr_selector2_31[1],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_497,addr_remain3_497);


wire[15:0] addr_selector3_498;
wire[15:0] addr_remain3_498;
address_decode_4 decoder_3_498 = address_decode_4(addr_selector2_31[2],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_498,addr_remain3_498);


wire[15:0] addr_selector3_499;
wire[15:0] addr_remain3_499;
address_decode_4 decoder_3_499 = address_decode_4(addr_selector2_31[3],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_499,addr_remain3_499);


wire[15:0] addr_selector3_500;
wire[15:0] addr_remain3_500;
address_decode_4 decoder_3_500 = address_decode_4(addr_selector2_31[4],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_500,addr_remain3_500);


wire[15:0] addr_selector3_501;
wire[15:0] addr_remain3_501;
address_decode_4 decoder_3_501 = address_decode_4(addr_selector2_31[5],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_501,addr_remain3_501);


wire[15:0] addr_selector3_502;
wire[15:0] addr_remain3_502;
address_decode_4 decoder_3_502 = address_decode_4(addr_selector2_31[6],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_502,addr_remain3_502);


wire[15:0] addr_selector3_503;
wire[15:0] addr_remain3_503;
address_decode_4 decoder_3_503 = address_decode_4(addr_selector2_31[7],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_503,addr_remain3_503);


wire[15:0] addr_selector3_504;
wire[15:0] addr_remain3_504;
address_decode_4 decoder_3_504 = address_decode_4(addr_selector2_31[8],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_504,addr_remain3_504);


wire[15:0] addr_selector3_505;
wire[15:0] addr_remain3_505;
address_decode_4 decoder_3_505 = address_decode_4(addr_selector2_31[9],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_505,addr_remain3_505);


wire[15:0] addr_selector3_506;
wire[15:0] addr_remain3_506;
address_decode_4 decoder_3_506 = address_decode_4(addr_selector2_31[10],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_506,addr_remain3_506);


wire[15:0] addr_selector3_507;
wire[15:0] addr_remain3_507;
address_decode_4 decoder_3_507 = address_decode_4(addr_selector2_31[11],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_507,addr_remain3_507);


wire[15:0] addr_selector3_508;
wire[15:0] addr_remain3_508;
address_decode_4 decoder_3_508 = address_decode_4(addr_selector2_31[12],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_508,addr_remain3_508);


wire[15:0] addr_selector3_509;
wire[15:0] addr_remain3_509;
address_decode_4 decoder_3_509 = address_decode_4(addr_selector2_31[13],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_509,addr_remain3_509);


wire[15:0] addr_selector3_510;
wire[15:0] addr_remain3_510;
address_decode_4 decoder_3_510 = address_decode_4(addr_selector2_31[14],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_510,addr_remain3_510);


wire[15:0] addr_selector3_511;
wire[15:0] addr_remain3_511;
address_decode_4 decoder_3_511 = address_decode_4(addr_selector2_31[15],addr_remain2_31[15:0],addr_remain2_31,addr_selector3_511,addr_remain3_511);


wire[15:0] addr_selector3_512;
wire[15:0] addr_remain3_512;
address_decode_4 decoder_3_512 = address_decode_4(addr_selector2_32[0],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_512,addr_remain3_512);


wire[15:0] addr_selector3_513;
wire[15:0] addr_remain3_513;
address_decode_4 decoder_3_513 = address_decode_4(addr_selector2_32[1],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_513,addr_remain3_513);


wire[15:0] addr_selector3_514;
wire[15:0] addr_remain3_514;
address_decode_4 decoder_3_514 = address_decode_4(addr_selector2_32[2],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_514,addr_remain3_514);


wire[15:0] addr_selector3_515;
wire[15:0] addr_remain3_515;
address_decode_4 decoder_3_515 = address_decode_4(addr_selector2_32[3],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_515,addr_remain3_515);


wire[15:0] addr_selector3_516;
wire[15:0] addr_remain3_516;
address_decode_4 decoder_3_516 = address_decode_4(addr_selector2_32[4],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_516,addr_remain3_516);


wire[15:0] addr_selector3_517;
wire[15:0] addr_remain3_517;
address_decode_4 decoder_3_517 = address_decode_4(addr_selector2_32[5],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_517,addr_remain3_517);


wire[15:0] addr_selector3_518;
wire[15:0] addr_remain3_518;
address_decode_4 decoder_3_518 = address_decode_4(addr_selector2_32[6],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_518,addr_remain3_518);


wire[15:0] addr_selector3_519;
wire[15:0] addr_remain3_519;
address_decode_4 decoder_3_519 = address_decode_4(addr_selector2_32[7],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_519,addr_remain3_519);


wire[15:0] addr_selector3_520;
wire[15:0] addr_remain3_520;
address_decode_4 decoder_3_520 = address_decode_4(addr_selector2_32[8],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_520,addr_remain3_520);


wire[15:0] addr_selector3_521;
wire[15:0] addr_remain3_521;
address_decode_4 decoder_3_521 = address_decode_4(addr_selector2_32[9],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_521,addr_remain3_521);


wire[15:0] addr_selector3_522;
wire[15:0] addr_remain3_522;
address_decode_4 decoder_3_522 = address_decode_4(addr_selector2_32[10],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_522,addr_remain3_522);


wire[15:0] addr_selector3_523;
wire[15:0] addr_remain3_523;
address_decode_4 decoder_3_523 = address_decode_4(addr_selector2_32[11],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_523,addr_remain3_523);


wire[15:0] addr_selector3_524;
wire[15:0] addr_remain3_524;
address_decode_4 decoder_3_524 = address_decode_4(addr_selector2_32[12],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_524,addr_remain3_524);


wire[15:0] addr_selector3_525;
wire[15:0] addr_remain3_525;
address_decode_4 decoder_3_525 = address_decode_4(addr_selector2_32[13],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_525,addr_remain3_525);


wire[15:0] addr_selector3_526;
wire[15:0] addr_remain3_526;
address_decode_4 decoder_3_526 = address_decode_4(addr_selector2_32[14],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_526,addr_remain3_526);


wire[15:0] addr_selector3_527;
wire[15:0] addr_remain3_527;
address_decode_4 decoder_3_527 = address_decode_4(addr_selector2_32[15],addr_remain2_32[15:0],addr_remain2_32,addr_selector3_527,addr_remain3_527);


wire[15:0] addr_selector3_528;
wire[15:0] addr_remain3_528;
address_decode_4 decoder_3_528 = address_decode_4(addr_selector2_33[0],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_528,addr_remain3_528);


wire[15:0] addr_selector3_529;
wire[15:0] addr_remain3_529;
address_decode_4 decoder_3_529 = address_decode_4(addr_selector2_33[1],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_529,addr_remain3_529);


wire[15:0] addr_selector3_530;
wire[15:0] addr_remain3_530;
address_decode_4 decoder_3_530 = address_decode_4(addr_selector2_33[2],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_530,addr_remain3_530);


wire[15:0] addr_selector3_531;
wire[15:0] addr_remain3_531;
address_decode_4 decoder_3_531 = address_decode_4(addr_selector2_33[3],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_531,addr_remain3_531);


wire[15:0] addr_selector3_532;
wire[15:0] addr_remain3_532;
address_decode_4 decoder_3_532 = address_decode_4(addr_selector2_33[4],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_532,addr_remain3_532);


wire[15:0] addr_selector3_533;
wire[15:0] addr_remain3_533;
address_decode_4 decoder_3_533 = address_decode_4(addr_selector2_33[5],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_533,addr_remain3_533);


wire[15:0] addr_selector3_534;
wire[15:0] addr_remain3_534;
address_decode_4 decoder_3_534 = address_decode_4(addr_selector2_33[6],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_534,addr_remain3_534);


wire[15:0] addr_selector3_535;
wire[15:0] addr_remain3_535;
address_decode_4 decoder_3_535 = address_decode_4(addr_selector2_33[7],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_535,addr_remain3_535);


wire[15:0] addr_selector3_536;
wire[15:0] addr_remain3_536;
address_decode_4 decoder_3_536 = address_decode_4(addr_selector2_33[8],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_536,addr_remain3_536);


wire[15:0] addr_selector3_537;
wire[15:0] addr_remain3_537;
address_decode_4 decoder_3_537 = address_decode_4(addr_selector2_33[9],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_537,addr_remain3_537);


wire[15:0] addr_selector3_538;
wire[15:0] addr_remain3_538;
address_decode_4 decoder_3_538 = address_decode_4(addr_selector2_33[10],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_538,addr_remain3_538);


wire[15:0] addr_selector3_539;
wire[15:0] addr_remain3_539;
address_decode_4 decoder_3_539 = address_decode_4(addr_selector2_33[11],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_539,addr_remain3_539);


wire[15:0] addr_selector3_540;
wire[15:0] addr_remain3_540;
address_decode_4 decoder_3_540 = address_decode_4(addr_selector2_33[12],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_540,addr_remain3_540);


wire[15:0] addr_selector3_541;
wire[15:0] addr_remain3_541;
address_decode_4 decoder_3_541 = address_decode_4(addr_selector2_33[13],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_541,addr_remain3_541);


wire[15:0] addr_selector3_542;
wire[15:0] addr_remain3_542;
address_decode_4 decoder_3_542 = address_decode_4(addr_selector2_33[14],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_542,addr_remain3_542);


wire[15:0] addr_selector3_543;
wire[15:0] addr_remain3_543;
address_decode_4 decoder_3_543 = address_decode_4(addr_selector2_33[15],addr_remain2_33[15:0],addr_remain2_33,addr_selector3_543,addr_remain3_543);


wire[15:0] addr_selector3_544;
wire[15:0] addr_remain3_544;
address_decode_4 decoder_3_544 = address_decode_4(addr_selector2_34[0],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_544,addr_remain3_544);


wire[15:0] addr_selector3_545;
wire[15:0] addr_remain3_545;
address_decode_4 decoder_3_545 = address_decode_4(addr_selector2_34[1],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_545,addr_remain3_545);


wire[15:0] addr_selector3_546;
wire[15:0] addr_remain3_546;
address_decode_4 decoder_3_546 = address_decode_4(addr_selector2_34[2],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_546,addr_remain3_546);


wire[15:0] addr_selector3_547;
wire[15:0] addr_remain3_547;
address_decode_4 decoder_3_547 = address_decode_4(addr_selector2_34[3],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_547,addr_remain3_547);


wire[15:0] addr_selector3_548;
wire[15:0] addr_remain3_548;
address_decode_4 decoder_3_548 = address_decode_4(addr_selector2_34[4],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_548,addr_remain3_548);


wire[15:0] addr_selector3_549;
wire[15:0] addr_remain3_549;
address_decode_4 decoder_3_549 = address_decode_4(addr_selector2_34[5],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_549,addr_remain3_549);


wire[15:0] addr_selector3_550;
wire[15:0] addr_remain3_550;
address_decode_4 decoder_3_550 = address_decode_4(addr_selector2_34[6],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_550,addr_remain3_550);


wire[15:0] addr_selector3_551;
wire[15:0] addr_remain3_551;
address_decode_4 decoder_3_551 = address_decode_4(addr_selector2_34[7],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_551,addr_remain3_551);


wire[15:0] addr_selector3_552;
wire[15:0] addr_remain3_552;
address_decode_4 decoder_3_552 = address_decode_4(addr_selector2_34[8],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_552,addr_remain3_552);


wire[15:0] addr_selector3_553;
wire[15:0] addr_remain3_553;
address_decode_4 decoder_3_553 = address_decode_4(addr_selector2_34[9],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_553,addr_remain3_553);


wire[15:0] addr_selector3_554;
wire[15:0] addr_remain3_554;
address_decode_4 decoder_3_554 = address_decode_4(addr_selector2_34[10],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_554,addr_remain3_554);


wire[15:0] addr_selector3_555;
wire[15:0] addr_remain3_555;
address_decode_4 decoder_3_555 = address_decode_4(addr_selector2_34[11],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_555,addr_remain3_555);


wire[15:0] addr_selector3_556;
wire[15:0] addr_remain3_556;
address_decode_4 decoder_3_556 = address_decode_4(addr_selector2_34[12],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_556,addr_remain3_556);


wire[15:0] addr_selector3_557;
wire[15:0] addr_remain3_557;
address_decode_4 decoder_3_557 = address_decode_4(addr_selector2_34[13],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_557,addr_remain3_557);


wire[15:0] addr_selector3_558;
wire[15:0] addr_remain3_558;
address_decode_4 decoder_3_558 = address_decode_4(addr_selector2_34[14],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_558,addr_remain3_558);


wire[15:0] addr_selector3_559;
wire[15:0] addr_remain3_559;
address_decode_4 decoder_3_559 = address_decode_4(addr_selector2_34[15],addr_remain2_34[15:0],addr_remain2_34,addr_selector3_559,addr_remain3_559);


wire[15:0] addr_selector3_560;
wire[15:0] addr_remain3_560;
address_decode_4 decoder_3_560 = address_decode_4(addr_selector2_35[0],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_560,addr_remain3_560);


wire[15:0] addr_selector3_561;
wire[15:0] addr_remain3_561;
address_decode_4 decoder_3_561 = address_decode_4(addr_selector2_35[1],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_561,addr_remain3_561);


wire[15:0] addr_selector3_562;
wire[15:0] addr_remain3_562;
address_decode_4 decoder_3_562 = address_decode_4(addr_selector2_35[2],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_562,addr_remain3_562);


wire[15:0] addr_selector3_563;
wire[15:0] addr_remain3_563;
address_decode_4 decoder_3_563 = address_decode_4(addr_selector2_35[3],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_563,addr_remain3_563);


wire[15:0] addr_selector3_564;
wire[15:0] addr_remain3_564;
address_decode_4 decoder_3_564 = address_decode_4(addr_selector2_35[4],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_564,addr_remain3_564);


wire[15:0] addr_selector3_565;
wire[15:0] addr_remain3_565;
address_decode_4 decoder_3_565 = address_decode_4(addr_selector2_35[5],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_565,addr_remain3_565);


wire[15:0] addr_selector3_566;
wire[15:0] addr_remain3_566;
address_decode_4 decoder_3_566 = address_decode_4(addr_selector2_35[6],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_566,addr_remain3_566);


wire[15:0] addr_selector3_567;
wire[15:0] addr_remain3_567;
address_decode_4 decoder_3_567 = address_decode_4(addr_selector2_35[7],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_567,addr_remain3_567);


wire[15:0] addr_selector3_568;
wire[15:0] addr_remain3_568;
address_decode_4 decoder_3_568 = address_decode_4(addr_selector2_35[8],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_568,addr_remain3_568);


wire[15:0] addr_selector3_569;
wire[15:0] addr_remain3_569;
address_decode_4 decoder_3_569 = address_decode_4(addr_selector2_35[9],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_569,addr_remain3_569);


wire[15:0] addr_selector3_570;
wire[15:0] addr_remain3_570;
address_decode_4 decoder_3_570 = address_decode_4(addr_selector2_35[10],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_570,addr_remain3_570);


wire[15:0] addr_selector3_571;
wire[15:0] addr_remain3_571;
address_decode_4 decoder_3_571 = address_decode_4(addr_selector2_35[11],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_571,addr_remain3_571);


wire[15:0] addr_selector3_572;
wire[15:0] addr_remain3_572;
address_decode_4 decoder_3_572 = address_decode_4(addr_selector2_35[12],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_572,addr_remain3_572);


wire[15:0] addr_selector3_573;
wire[15:0] addr_remain3_573;
address_decode_4 decoder_3_573 = address_decode_4(addr_selector2_35[13],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_573,addr_remain3_573);


wire[15:0] addr_selector3_574;
wire[15:0] addr_remain3_574;
address_decode_4 decoder_3_574 = address_decode_4(addr_selector2_35[14],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_574,addr_remain3_574);


wire[15:0] addr_selector3_575;
wire[15:0] addr_remain3_575;
address_decode_4 decoder_3_575 = address_decode_4(addr_selector2_35[15],addr_remain2_35[15:0],addr_remain2_35,addr_selector3_575,addr_remain3_575);


wire[15:0] addr_selector3_576;
wire[15:0] addr_remain3_576;
address_decode_4 decoder_3_576 = address_decode_4(addr_selector2_36[0],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_576,addr_remain3_576);


wire[15:0] addr_selector3_577;
wire[15:0] addr_remain3_577;
address_decode_4 decoder_3_577 = address_decode_4(addr_selector2_36[1],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_577,addr_remain3_577);


wire[15:0] addr_selector3_578;
wire[15:0] addr_remain3_578;
address_decode_4 decoder_3_578 = address_decode_4(addr_selector2_36[2],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_578,addr_remain3_578);


wire[15:0] addr_selector3_579;
wire[15:0] addr_remain3_579;
address_decode_4 decoder_3_579 = address_decode_4(addr_selector2_36[3],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_579,addr_remain3_579);


wire[15:0] addr_selector3_580;
wire[15:0] addr_remain3_580;
address_decode_4 decoder_3_580 = address_decode_4(addr_selector2_36[4],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_580,addr_remain3_580);


wire[15:0] addr_selector3_581;
wire[15:0] addr_remain3_581;
address_decode_4 decoder_3_581 = address_decode_4(addr_selector2_36[5],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_581,addr_remain3_581);


wire[15:0] addr_selector3_582;
wire[15:0] addr_remain3_582;
address_decode_4 decoder_3_582 = address_decode_4(addr_selector2_36[6],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_582,addr_remain3_582);


wire[15:0] addr_selector3_583;
wire[15:0] addr_remain3_583;
address_decode_4 decoder_3_583 = address_decode_4(addr_selector2_36[7],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_583,addr_remain3_583);


wire[15:0] addr_selector3_584;
wire[15:0] addr_remain3_584;
address_decode_4 decoder_3_584 = address_decode_4(addr_selector2_36[8],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_584,addr_remain3_584);


wire[15:0] addr_selector3_585;
wire[15:0] addr_remain3_585;
address_decode_4 decoder_3_585 = address_decode_4(addr_selector2_36[9],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_585,addr_remain3_585);


wire[15:0] addr_selector3_586;
wire[15:0] addr_remain3_586;
address_decode_4 decoder_3_586 = address_decode_4(addr_selector2_36[10],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_586,addr_remain3_586);


wire[15:0] addr_selector3_587;
wire[15:0] addr_remain3_587;
address_decode_4 decoder_3_587 = address_decode_4(addr_selector2_36[11],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_587,addr_remain3_587);


wire[15:0] addr_selector3_588;
wire[15:0] addr_remain3_588;
address_decode_4 decoder_3_588 = address_decode_4(addr_selector2_36[12],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_588,addr_remain3_588);


wire[15:0] addr_selector3_589;
wire[15:0] addr_remain3_589;
address_decode_4 decoder_3_589 = address_decode_4(addr_selector2_36[13],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_589,addr_remain3_589);


wire[15:0] addr_selector3_590;
wire[15:0] addr_remain3_590;
address_decode_4 decoder_3_590 = address_decode_4(addr_selector2_36[14],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_590,addr_remain3_590);


wire[15:0] addr_selector3_591;
wire[15:0] addr_remain3_591;
address_decode_4 decoder_3_591 = address_decode_4(addr_selector2_36[15],addr_remain2_36[15:0],addr_remain2_36,addr_selector3_591,addr_remain3_591);


wire[15:0] addr_selector3_592;
wire[15:0] addr_remain3_592;
address_decode_4 decoder_3_592 = address_decode_4(addr_selector2_37[0],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_592,addr_remain3_592);


wire[15:0] addr_selector3_593;
wire[15:0] addr_remain3_593;
address_decode_4 decoder_3_593 = address_decode_4(addr_selector2_37[1],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_593,addr_remain3_593);


wire[15:0] addr_selector3_594;
wire[15:0] addr_remain3_594;
address_decode_4 decoder_3_594 = address_decode_4(addr_selector2_37[2],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_594,addr_remain3_594);


wire[15:0] addr_selector3_595;
wire[15:0] addr_remain3_595;
address_decode_4 decoder_3_595 = address_decode_4(addr_selector2_37[3],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_595,addr_remain3_595);


wire[15:0] addr_selector3_596;
wire[15:0] addr_remain3_596;
address_decode_4 decoder_3_596 = address_decode_4(addr_selector2_37[4],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_596,addr_remain3_596);


wire[15:0] addr_selector3_597;
wire[15:0] addr_remain3_597;
address_decode_4 decoder_3_597 = address_decode_4(addr_selector2_37[5],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_597,addr_remain3_597);


wire[15:0] addr_selector3_598;
wire[15:0] addr_remain3_598;
address_decode_4 decoder_3_598 = address_decode_4(addr_selector2_37[6],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_598,addr_remain3_598);


wire[15:0] addr_selector3_599;
wire[15:0] addr_remain3_599;
address_decode_4 decoder_3_599 = address_decode_4(addr_selector2_37[7],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_599,addr_remain3_599);


wire[15:0] addr_selector3_600;
wire[15:0] addr_remain3_600;
address_decode_4 decoder_3_600 = address_decode_4(addr_selector2_37[8],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_600,addr_remain3_600);


wire[15:0] addr_selector3_601;
wire[15:0] addr_remain3_601;
address_decode_4 decoder_3_601 = address_decode_4(addr_selector2_37[9],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_601,addr_remain3_601);


wire[15:0] addr_selector3_602;
wire[15:0] addr_remain3_602;
address_decode_4 decoder_3_602 = address_decode_4(addr_selector2_37[10],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_602,addr_remain3_602);


wire[15:0] addr_selector3_603;
wire[15:0] addr_remain3_603;
address_decode_4 decoder_3_603 = address_decode_4(addr_selector2_37[11],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_603,addr_remain3_603);


wire[15:0] addr_selector3_604;
wire[15:0] addr_remain3_604;
address_decode_4 decoder_3_604 = address_decode_4(addr_selector2_37[12],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_604,addr_remain3_604);


wire[15:0] addr_selector3_605;
wire[15:0] addr_remain3_605;
address_decode_4 decoder_3_605 = address_decode_4(addr_selector2_37[13],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_605,addr_remain3_605);


wire[15:0] addr_selector3_606;
wire[15:0] addr_remain3_606;
address_decode_4 decoder_3_606 = address_decode_4(addr_selector2_37[14],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_606,addr_remain3_606);


wire[15:0] addr_selector3_607;
wire[15:0] addr_remain3_607;
address_decode_4 decoder_3_607 = address_decode_4(addr_selector2_37[15],addr_remain2_37[15:0],addr_remain2_37,addr_selector3_607,addr_remain3_607);


wire[15:0] addr_selector3_608;
wire[15:0] addr_remain3_608;
address_decode_4 decoder_3_608 = address_decode_4(addr_selector2_38[0],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_608,addr_remain3_608);


wire[15:0] addr_selector3_609;
wire[15:0] addr_remain3_609;
address_decode_4 decoder_3_609 = address_decode_4(addr_selector2_38[1],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_609,addr_remain3_609);


wire[15:0] addr_selector3_610;
wire[15:0] addr_remain3_610;
address_decode_4 decoder_3_610 = address_decode_4(addr_selector2_38[2],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_610,addr_remain3_610);


wire[15:0] addr_selector3_611;
wire[15:0] addr_remain3_611;
address_decode_4 decoder_3_611 = address_decode_4(addr_selector2_38[3],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_611,addr_remain3_611);


wire[15:0] addr_selector3_612;
wire[15:0] addr_remain3_612;
address_decode_4 decoder_3_612 = address_decode_4(addr_selector2_38[4],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_612,addr_remain3_612);


wire[15:0] addr_selector3_613;
wire[15:0] addr_remain3_613;
address_decode_4 decoder_3_613 = address_decode_4(addr_selector2_38[5],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_613,addr_remain3_613);


wire[15:0] addr_selector3_614;
wire[15:0] addr_remain3_614;
address_decode_4 decoder_3_614 = address_decode_4(addr_selector2_38[6],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_614,addr_remain3_614);


wire[15:0] addr_selector3_615;
wire[15:0] addr_remain3_615;
address_decode_4 decoder_3_615 = address_decode_4(addr_selector2_38[7],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_615,addr_remain3_615);


wire[15:0] addr_selector3_616;
wire[15:0] addr_remain3_616;
address_decode_4 decoder_3_616 = address_decode_4(addr_selector2_38[8],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_616,addr_remain3_616);


wire[15:0] addr_selector3_617;
wire[15:0] addr_remain3_617;
address_decode_4 decoder_3_617 = address_decode_4(addr_selector2_38[9],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_617,addr_remain3_617);


wire[15:0] addr_selector3_618;
wire[15:0] addr_remain3_618;
address_decode_4 decoder_3_618 = address_decode_4(addr_selector2_38[10],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_618,addr_remain3_618);


wire[15:0] addr_selector3_619;
wire[15:0] addr_remain3_619;
address_decode_4 decoder_3_619 = address_decode_4(addr_selector2_38[11],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_619,addr_remain3_619);


wire[15:0] addr_selector3_620;
wire[15:0] addr_remain3_620;
address_decode_4 decoder_3_620 = address_decode_4(addr_selector2_38[12],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_620,addr_remain3_620);


wire[15:0] addr_selector3_621;
wire[15:0] addr_remain3_621;
address_decode_4 decoder_3_621 = address_decode_4(addr_selector2_38[13],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_621,addr_remain3_621);


wire[15:0] addr_selector3_622;
wire[15:0] addr_remain3_622;
address_decode_4 decoder_3_622 = address_decode_4(addr_selector2_38[14],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_622,addr_remain3_622);


wire[15:0] addr_selector3_623;
wire[15:0] addr_remain3_623;
address_decode_4 decoder_3_623 = address_decode_4(addr_selector2_38[15],addr_remain2_38[15:0],addr_remain2_38,addr_selector3_623,addr_remain3_623);


wire[15:0] addr_selector3_624;
wire[15:0] addr_remain3_624;
address_decode_4 decoder_3_624 = address_decode_4(addr_selector2_39[0],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_624,addr_remain3_624);


wire[15:0] addr_selector3_625;
wire[15:0] addr_remain3_625;
address_decode_4 decoder_3_625 = address_decode_4(addr_selector2_39[1],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_625,addr_remain3_625);


wire[15:0] addr_selector3_626;
wire[15:0] addr_remain3_626;
address_decode_4 decoder_3_626 = address_decode_4(addr_selector2_39[2],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_626,addr_remain3_626);


wire[15:0] addr_selector3_627;
wire[15:0] addr_remain3_627;
address_decode_4 decoder_3_627 = address_decode_4(addr_selector2_39[3],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_627,addr_remain3_627);


wire[15:0] addr_selector3_628;
wire[15:0] addr_remain3_628;
address_decode_4 decoder_3_628 = address_decode_4(addr_selector2_39[4],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_628,addr_remain3_628);


wire[15:0] addr_selector3_629;
wire[15:0] addr_remain3_629;
address_decode_4 decoder_3_629 = address_decode_4(addr_selector2_39[5],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_629,addr_remain3_629);


wire[15:0] addr_selector3_630;
wire[15:0] addr_remain3_630;
address_decode_4 decoder_3_630 = address_decode_4(addr_selector2_39[6],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_630,addr_remain3_630);


wire[15:0] addr_selector3_631;
wire[15:0] addr_remain3_631;
address_decode_4 decoder_3_631 = address_decode_4(addr_selector2_39[7],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_631,addr_remain3_631);


wire[15:0] addr_selector3_632;
wire[15:0] addr_remain3_632;
address_decode_4 decoder_3_632 = address_decode_4(addr_selector2_39[8],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_632,addr_remain3_632);


wire[15:0] addr_selector3_633;
wire[15:0] addr_remain3_633;
address_decode_4 decoder_3_633 = address_decode_4(addr_selector2_39[9],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_633,addr_remain3_633);


wire[15:0] addr_selector3_634;
wire[15:0] addr_remain3_634;
address_decode_4 decoder_3_634 = address_decode_4(addr_selector2_39[10],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_634,addr_remain3_634);


wire[15:0] addr_selector3_635;
wire[15:0] addr_remain3_635;
address_decode_4 decoder_3_635 = address_decode_4(addr_selector2_39[11],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_635,addr_remain3_635);


wire[15:0] addr_selector3_636;
wire[15:0] addr_remain3_636;
address_decode_4 decoder_3_636 = address_decode_4(addr_selector2_39[12],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_636,addr_remain3_636);


wire[15:0] addr_selector3_637;
wire[15:0] addr_remain3_637;
address_decode_4 decoder_3_637 = address_decode_4(addr_selector2_39[13],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_637,addr_remain3_637);


wire[15:0] addr_selector3_638;
wire[15:0] addr_remain3_638;
address_decode_4 decoder_3_638 = address_decode_4(addr_selector2_39[14],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_638,addr_remain3_638);


wire[15:0] addr_selector3_639;
wire[15:0] addr_remain3_639;
address_decode_4 decoder_3_639 = address_decode_4(addr_selector2_39[15],addr_remain2_39[15:0],addr_remain2_39,addr_selector3_639,addr_remain3_639);


wire[15:0] addr_selector3_640;
wire[15:0] addr_remain3_640;
address_decode_4 decoder_3_640 = address_decode_4(addr_selector2_40[0],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_640,addr_remain3_640);


wire[15:0] addr_selector3_641;
wire[15:0] addr_remain3_641;
address_decode_4 decoder_3_641 = address_decode_4(addr_selector2_40[1],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_641,addr_remain3_641);


wire[15:0] addr_selector3_642;
wire[15:0] addr_remain3_642;
address_decode_4 decoder_3_642 = address_decode_4(addr_selector2_40[2],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_642,addr_remain3_642);


wire[15:0] addr_selector3_643;
wire[15:0] addr_remain3_643;
address_decode_4 decoder_3_643 = address_decode_4(addr_selector2_40[3],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_643,addr_remain3_643);


wire[15:0] addr_selector3_644;
wire[15:0] addr_remain3_644;
address_decode_4 decoder_3_644 = address_decode_4(addr_selector2_40[4],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_644,addr_remain3_644);


wire[15:0] addr_selector3_645;
wire[15:0] addr_remain3_645;
address_decode_4 decoder_3_645 = address_decode_4(addr_selector2_40[5],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_645,addr_remain3_645);


wire[15:0] addr_selector3_646;
wire[15:0] addr_remain3_646;
address_decode_4 decoder_3_646 = address_decode_4(addr_selector2_40[6],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_646,addr_remain3_646);


wire[15:0] addr_selector3_647;
wire[15:0] addr_remain3_647;
address_decode_4 decoder_3_647 = address_decode_4(addr_selector2_40[7],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_647,addr_remain3_647);


wire[15:0] addr_selector3_648;
wire[15:0] addr_remain3_648;
address_decode_4 decoder_3_648 = address_decode_4(addr_selector2_40[8],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_648,addr_remain3_648);


wire[15:0] addr_selector3_649;
wire[15:0] addr_remain3_649;
address_decode_4 decoder_3_649 = address_decode_4(addr_selector2_40[9],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_649,addr_remain3_649);


wire[15:0] addr_selector3_650;
wire[15:0] addr_remain3_650;
address_decode_4 decoder_3_650 = address_decode_4(addr_selector2_40[10],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_650,addr_remain3_650);


wire[15:0] addr_selector3_651;
wire[15:0] addr_remain3_651;
address_decode_4 decoder_3_651 = address_decode_4(addr_selector2_40[11],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_651,addr_remain3_651);


wire[15:0] addr_selector3_652;
wire[15:0] addr_remain3_652;
address_decode_4 decoder_3_652 = address_decode_4(addr_selector2_40[12],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_652,addr_remain3_652);


wire[15:0] addr_selector3_653;
wire[15:0] addr_remain3_653;
address_decode_4 decoder_3_653 = address_decode_4(addr_selector2_40[13],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_653,addr_remain3_653);


wire[15:0] addr_selector3_654;
wire[15:0] addr_remain3_654;
address_decode_4 decoder_3_654 = address_decode_4(addr_selector2_40[14],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_654,addr_remain3_654);


wire[15:0] addr_selector3_655;
wire[15:0] addr_remain3_655;
address_decode_4 decoder_3_655 = address_decode_4(addr_selector2_40[15],addr_remain2_40[15:0],addr_remain2_40,addr_selector3_655,addr_remain3_655);


wire[15:0] addr_selector3_656;
wire[15:0] addr_remain3_656;
address_decode_4 decoder_3_656 = address_decode_4(addr_selector2_41[0],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_656,addr_remain3_656);


wire[15:0] addr_selector3_657;
wire[15:0] addr_remain3_657;
address_decode_4 decoder_3_657 = address_decode_4(addr_selector2_41[1],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_657,addr_remain3_657);


wire[15:0] addr_selector3_658;
wire[15:0] addr_remain3_658;
address_decode_4 decoder_3_658 = address_decode_4(addr_selector2_41[2],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_658,addr_remain3_658);


wire[15:0] addr_selector3_659;
wire[15:0] addr_remain3_659;
address_decode_4 decoder_3_659 = address_decode_4(addr_selector2_41[3],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_659,addr_remain3_659);


wire[15:0] addr_selector3_660;
wire[15:0] addr_remain3_660;
address_decode_4 decoder_3_660 = address_decode_4(addr_selector2_41[4],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_660,addr_remain3_660);


wire[15:0] addr_selector3_661;
wire[15:0] addr_remain3_661;
address_decode_4 decoder_3_661 = address_decode_4(addr_selector2_41[5],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_661,addr_remain3_661);


wire[15:0] addr_selector3_662;
wire[15:0] addr_remain3_662;
address_decode_4 decoder_3_662 = address_decode_4(addr_selector2_41[6],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_662,addr_remain3_662);


wire[15:0] addr_selector3_663;
wire[15:0] addr_remain3_663;
address_decode_4 decoder_3_663 = address_decode_4(addr_selector2_41[7],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_663,addr_remain3_663);


wire[15:0] addr_selector3_664;
wire[15:0] addr_remain3_664;
address_decode_4 decoder_3_664 = address_decode_4(addr_selector2_41[8],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_664,addr_remain3_664);


wire[15:0] addr_selector3_665;
wire[15:0] addr_remain3_665;
address_decode_4 decoder_3_665 = address_decode_4(addr_selector2_41[9],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_665,addr_remain3_665);


wire[15:0] addr_selector3_666;
wire[15:0] addr_remain3_666;
address_decode_4 decoder_3_666 = address_decode_4(addr_selector2_41[10],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_666,addr_remain3_666);


wire[15:0] addr_selector3_667;
wire[15:0] addr_remain3_667;
address_decode_4 decoder_3_667 = address_decode_4(addr_selector2_41[11],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_667,addr_remain3_667);


wire[15:0] addr_selector3_668;
wire[15:0] addr_remain3_668;
address_decode_4 decoder_3_668 = address_decode_4(addr_selector2_41[12],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_668,addr_remain3_668);


wire[15:0] addr_selector3_669;
wire[15:0] addr_remain3_669;
address_decode_4 decoder_3_669 = address_decode_4(addr_selector2_41[13],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_669,addr_remain3_669);


wire[15:0] addr_selector3_670;
wire[15:0] addr_remain3_670;
address_decode_4 decoder_3_670 = address_decode_4(addr_selector2_41[14],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_670,addr_remain3_670);


wire[15:0] addr_selector3_671;
wire[15:0] addr_remain3_671;
address_decode_4 decoder_3_671 = address_decode_4(addr_selector2_41[15],addr_remain2_41[15:0],addr_remain2_41,addr_selector3_671,addr_remain3_671);


wire[15:0] addr_selector3_672;
wire[15:0] addr_remain3_672;
address_decode_4 decoder_3_672 = address_decode_4(addr_selector2_42[0],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_672,addr_remain3_672);


wire[15:0] addr_selector3_673;
wire[15:0] addr_remain3_673;
address_decode_4 decoder_3_673 = address_decode_4(addr_selector2_42[1],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_673,addr_remain3_673);


wire[15:0] addr_selector3_674;
wire[15:0] addr_remain3_674;
address_decode_4 decoder_3_674 = address_decode_4(addr_selector2_42[2],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_674,addr_remain3_674);


wire[15:0] addr_selector3_675;
wire[15:0] addr_remain3_675;
address_decode_4 decoder_3_675 = address_decode_4(addr_selector2_42[3],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_675,addr_remain3_675);


wire[15:0] addr_selector3_676;
wire[15:0] addr_remain3_676;
address_decode_4 decoder_3_676 = address_decode_4(addr_selector2_42[4],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_676,addr_remain3_676);


wire[15:0] addr_selector3_677;
wire[15:0] addr_remain3_677;
address_decode_4 decoder_3_677 = address_decode_4(addr_selector2_42[5],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_677,addr_remain3_677);


wire[15:0] addr_selector3_678;
wire[15:0] addr_remain3_678;
address_decode_4 decoder_3_678 = address_decode_4(addr_selector2_42[6],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_678,addr_remain3_678);


wire[15:0] addr_selector3_679;
wire[15:0] addr_remain3_679;
address_decode_4 decoder_3_679 = address_decode_4(addr_selector2_42[7],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_679,addr_remain3_679);


wire[15:0] addr_selector3_680;
wire[15:0] addr_remain3_680;
address_decode_4 decoder_3_680 = address_decode_4(addr_selector2_42[8],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_680,addr_remain3_680);


wire[15:0] addr_selector3_681;
wire[15:0] addr_remain3_681;
address_decode_4 decoder_3_681 = address_decode_4(addr_selector2_42[9],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_681,addr_remain3_681);


wire[15:0] addr_selector3_682;
wire[15:0] addr_remain3_682;
address_decode_4 decoder_3_682 = address_decode_4(addr_selector2_42[10],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_682,addr_remain3_682);


wire[15:0] addr_selector3_683;
wire[15:0] addr_remain3_683;
address_decode_4 decoder_3_683 = address_decode_4(addr_selector2_42[11],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_683,addr_remain3_683);


wire[15:0] addr_selector3_684;
wire[15:0] addr_remain3_684;
address_decode_4 decoder_3_684 = address_decode_4(addr_selector2_42[12],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_684,addr_remain3_684);


wire[15:0] addr_selector3_685;
wire[15:0] addr_remain3_685;
address_decode_4 decoder_3_685 = address_decode_4(addr_selector2_42[13],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_685,addr_remain3_685);


wire[15:0] addr_selector3_686;
wire[15:0] addr_remain3_686;
address_decode_4 decoder_3_686 = address_decode_4(addr_selector2_42[14],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_686,addr_remain3_686);


wire[15:0] addr_selector3_687;
wire[15:0] addr_remain3_687;
address_decode_4 decoder_3_687 = address_decode_4(addr_selector2_42[15],addr_remain2_42[15:0],addr_remain2_42,addr_selector3_687,addr_remain3_687);


wire[15:0] addr_selector3_688;
wire[15:0] addr_remain3_688;
address_decode_4 decoder_3_688 = address_decode_4(addr_selector2_43[0],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_688,addr_remain3_688);


wire[15:0] addr_selector3_689;
wire[15:0] addr_remain3_689;
address_decode_4 decoder_3_689 = address_decode_4(addr_selector2_43[1],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_689,addr_remain3_689);


wire[15:0] addr_selector3_690;
wire[15:0] addr_remain3_690;
address_decode_4 decoder_3_690 = address_decode_4(addr_selector2_43[2],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_690,addr_remain3_690);


wire[15:0] addr_selector3_691;
wire[15:0] addr_remain3_691;
address_decode_4 decoder_3_691 = address_decode_4(addr_selector2_43[3],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_691,addr_remain3_691);


wire[15:0] addr_selector3_692;
wire[15:0] addr_remain3_692;
address_decode_4 decoder_3_692 = address_decode_4(addr_selector2_43[4],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_692,addr_remain3_692);


wire[15:0] addr_selector3_693;
wire[15:0] addr_remain3_693;
address_decode_4 decoder_3_693 = address_decode_4(addr_selector2_43[5],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_693,addr_remain3_693);


wire[15:0] addr_selector3_694;
wire[15:0] addr_remain3_694;
address_decode_4 decoder_3_694 = address_decode_4(addr_selector2_43[6],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_694,addr_remain3_694);


wire[15:0] addr_selector3_695;
wire[15:0] addr_remain3_695;
address_decode_4 decoder_3_695 = address_decode_4(addr_selector2_43[7],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_695,addr_remain3_695);


wire[15:0] addr_selector3_696;
wire[15:0] addr_remain3_696;
address_decode_4 decoder_3_696 = address_decode_4(addr_selector2_43[8],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_696,addr_remain3_696);


wire[15:0] addr_selector3_697;
wire[15:0] addr_remain3_697;
address_decode_4 decoder_3_697 = address_decode_4(addr_selector2_43[9],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_697,addr_remain3_697);


wire[15:0] addr_selector3_698;
wire[15:0] addr_remain3_698;
address_decode_4 decoder_3_698 = address_decode_4(addr_selector2_43[10],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_698,addr_remain3_698);


wire[15:0] addr_selector3_699;
wire[15:0] addr_remain3_699;
address_decode_4 decoder_3_699 = address_decode_4(addr_selector2_43[11],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_699,addr_remain3_699);


wire[15:0] addr_selector3_700;
wire[15:0] addr_remain3_700;
address_decode_4 decoder_3_700 = address_decode_4(addr_selector2_43[12],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_700,addr_remain3_700);


wire[15:0] addr_selector3_701;
wire[15:0] addr_remain3_701;
address_decode_4 decoder_3_701 = address_decode_4(addr_selector2_43[13],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_701,addr_remain3_701);


wire[15:0] addr_selector3_702;
wire[15:0] addr_remain3_702;
address_decode_4 decoder_3_702 = address_decode_4(addr_selector2_43[14],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_702,addr_remain3_702);


wire[15:0] addr_selector3_703;
wire[15:0] addr_remain3_703;
address_decode_4 decoder_3_703 = address_decode_4(addr_selector2_43[15],addr_remain2_43[15:0],addr_remain2_43,addr_selector3_703,addr_remain3_703);


wire[15:0] addr_selector3_704;
wire[15:0] addr_remain3_704;
address_decode_4 decoder_3_704 = address_decode_4(addr_selector2_44[0],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_704,addr_remain3_704);


wire[15:0] addr_selector3_705;
wire[15:0] addr_remain3_705;
address_decode_4 decoder_3_705 = address_decode_4(addr_selector2_44[1],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_705,addr_remain3_705);


wire[15:0] addr_selector3_706;
wire[15:0] addr_remain3_706;
address_decode_4 decoder_3_706 = address_decode_4(addr_selector2_44[2],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_706,addr_remain3_706);


wire[15:0] addr_selector3_707;
wire[15:0] addr_remain3_707;
address_decode_4 decoder_3_707 = address_decode_4(addr_selector2_44[3],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_707,addr_remain3_707);


wire[15:0] addr_selector3_708;
wire[15:0] addr_remain3_708;
address_decode_4 decoder_3_708 = address_decode_4(addr_selector2_44[4],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_708,addr_remain3_708);


wire[15:0] addr_selector3_709;
wire[15:0] addr_remain3_709;
address_decode_4 decoder_3_709 = address_decode_4(addr_selector2_44[5],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_709,addr_remain3_709);


wire[15:0] addr_selector3_710;
wire[15:0] addr_remain3_710;
address_decode_4 decoder_3_710 = address_decode_4(addr_selector2_44[6],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_710,addr_remain3_710);


wire[15:0] addr_selector3_711;
wire[15:0] addr_remain3_711;
address_decode_4 decoder_3_711 = address_decode_4(addr_selector2_44[7],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_711,addr_remain3_711);


wire[15:0] addr_selector3_712;
wire[15:0] addr_remain3_712;
address_decode_4 decoder_3_712 = address_decode_4(addr_selector2_44[8],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_712,addr_remain3_712);


wire[15:0] addr_selector3_713;
wire[15:0] addr_remain3_713;
address_decode_4 decoder_3_713 = address_decode_4(addr_selector2_44[9],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_713,addr_remain3_713);


wire[15:0] addr_selector3_714;
wire[15:0] addr_remain3_714;
address_decode_4 decoder_3_714 = address_decode_4(addr_selector2_44[10],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_714,addr_remain3_714);


wire[15:0] addr_selector3_715;
wire[15:0] addr_remain3_715;
address_decode_4 decoder_3_715 = address_decode_4(addr_selector2_44[11],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_715,addr_remain3_715);


wire[15:0] addr_selector3_716;
wire[15:0] addr_remain3_716;
address_decode_4 decoder_3_716 = address_decode_4(addr_selector2_44[12],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_716,addr_remain3_716);


wire[15:0] addr_selector3_717;
wire[15:0] addr_remain3_717;
address_decode_4 decoder_3_717 = address_decode_4(addr_selector2_44[13],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_717,addr_remain3_717);


wire[15:0] addr_selector3_718;
wire[15:0] addr_remain3_718;
address_decode_4 decoder_3_718 = address_decode_4(addr_selector2_44[14],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_718,addr_remain3_718);


wire[15:0] addr_selector3_719;
wire[15:0] addr_remain3_719;
address_decode_4 decoder_3_719 = address_decode_4(addr_selector2_44[15],addr_remain2_44[15:0],addr_remain2_44,addr_selector3_719,addr_remain3_719);


wire[15:0] addr_selector3_720;
wire[15:0] addr_remain3_720;
address_decode_4 decoder_3_720 = address_decode_4(addr_selector2_45[0],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_720,addr_remain3_720);


wire[15:0] addr_selector3_721;
wire[15:0] addr_remain3_721;
address_decode_4 decoder_3_721 = address_decode_4(addr_selector2_45[1],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_721,addr_remain3_721);


wire[15:0] addr_selector3_722;
wire[15:0] addr_remain3_722;
address_decode_4 decoder_3_722 = address_decode_4(addr_selector2_45[2],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_722,addr_remain3_722);


wire[15:0] addr_selector3_723;
wire[15:0] addr_remain3_723;
address_decode_4 decoder_3_723 = address_decode_4(addr_selector2_45[3],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_723,addr_remain3_723);


wire[15:0] addr_selector3_724;
wire[15:0] addr_remain3_724;
address_decode_4 decoder_3_724 = address_decode_4(addr_selector2_45[4],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_724,addr_remain3_724);


wire[15:0] addr_selector3_725;
wire[15:0] addr_remain3_725;
address_decode_4 decoder_3_725 = address_decode_4(addr_selector2_45[5],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_725,addr_remain3_725);


wire[15:0] addr_selector3_726;
wire[15:0] addr_remain3_726;
address_decode_4 decoder_3_726 = address_decode_4(addr_selector2_45[6],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_726,addr_remain3_726);


wire[15:0] addr_selector3_727;
wire[15:0] addr_remain3_727;
address_decode_4 decoder_3_727 = address_decode_4(addr_selector2_45[7],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_727,addr_remain3_727);


wire[15:0] addr_selector3_728;
wire[15:0] addr_remain3_728;
address_decode_4 decoder_3_728 = address_decode_4(addr_selector2_45[8],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_728,addr_remain3_728);


wire[15:0] addr_selector3_729;
wire[15:0] addr_remain3_729;
address_decode_4 decoder_3_729 = address_decode_4(addr_selector2_45[9],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_729,addr_remain3_729);


wire[15:0] addr_selector3_730;
wire[15:0] addr_remain3_730;
address_decode_4 decoder_3_730 = address_decode_4(addr_selector2_45[10],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_730,addr_remain3_730);


wire[15:0] addr_selector3_731;
wire[15:0] addr_remain3_731;
address_decode_4 decoder_3_731 = address_decode_4(addr_selector2_45[11],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_731,addr_remain3_731);


wire[15:0] addr_selector3_732;
wire[15:0] addr_remain3_732;
address_decode_4 decoder_3_732 = address_decode_4(addr_selector2_45[12],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_732,addr_remain3_732);


wire[15:0] addr_selector3_733;
wire[15:0] addr_remain3_733;
address_decode_4 decoder_3_733 = address_decode_4(addr_selector2_45[13],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_733,addr_remain3_733);


wire[15:0] addr_selector3_734;
wire[15:0] addr_remain3_734;
address_decode_4 decoder_3_734 = address_decode_4(addr_selector2_45[14],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_734,addr_remain3_734);


wire[15:0] addr_selector3_735;
wire[15:0] addr_remain3_735;
address_decode_4 decoder_3_735 = address_decode_4(addr_selector2_45[15],addr_remain2_45[15:0],addr_remain2_45,addr_selector3_735,addr_remain3_735);


wire[15:0] addr_selector3_736;
wire[15:0] addr_remain3_736;
address_decode_4 decoder_3_736 = address_decode_4(addr_selector2_46[0],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_736,addr_remain3_736);


wire[15:0] addr_selector3_737;
wire[15:0] addr_remain3_737;
address_decode_4 decoder_3_737 = address_decode_4(addr_selector2_46[1],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_737,addr_remain3_737);


wire[15:0] addr_selector3_738;
wire[15:0] addr_remain3_738;
address_decode_4 decoder_3_738 = address_decode_4(addr_selector2_46[2],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_738,addr_remain3_738);


wire[15:0] addr_selector3_739;
wire[15:0] addr_remain3_739;
address_decode_4 decoder_3_739 = address_decode_4(addr_selector2_46[3],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_739,addr_remain3_739);


wire[15:0] addr_selector3_740;
wire[15:0] addr_remain3_740;
address_decode_4 decoder_3_740 = address_decode_4(addr_selector2_46[4],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_740,addr_remain3_740);


wire[15:0] addr_selector3_741;
wire[15:0] addr_remain3_741;
address_decode_4 decoder_3_741 = address_decode_4(addr_selector2_46[5],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_741,addr_remain3_741);


wire[15:0] addr_selector3_742;
wire[15:0] addr_remain3_742;
address_decode_4 decoder_3_742 = address_decode_4(addr_selector2_46[6],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_742,addr_remain3_742);


wire[15:0] addr_selector3_743;
wire[15:0] addr_remain3_743;
address_decode_4 decoder_3_743 = address_decode_4(addr_selector2_46[7],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_743,addr_remain3_743);


wire[15:0] addr_selector3_744;
wire[15:0] addr_remain3_744;
address_decode_4 decoder_3_744 = address_decode_4(addr_selector2_46[8],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_744,addr_remain3_744);


wire[15:0] addr_selector3_745;
wire[15:0] addr_remain3_745;
address_decode_4 decoder_3_745 = address_decode_4(addr_selector2_46[9],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_745,addr_remain3_745);


wire[15:0] addr_selector3_746;
wire[15:0] addr_remain3_746;
address_decode_4 decoder_3_746 = address_decode_4(addr_selector2_46[10],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_746,addr_remain3_746);


wire[15:0] addr_selector3_747;
wire[15:0] addr_remain3_747;
address_decode_4 decoder_3_747 = address_decode_4(addr_selector2_46[11],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_747,addr_remain3_747);


wire[15:0] addr_selector3_748;
wire[15:0] addr_remain3_748;
address_decode_4 decoder_3_748 = address_decode_4(addr_selector2_46[12],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_748,addr_remain3_748);


wire[15:0] addr_selector3_749;
wire[15:0] addr_remain3_749;
address_decode_4 decoder_3_749 = address_decode_4(addr_selector2_46[13],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_749,addr_remain3_749);


wire[15:0] addr_selector3_750;
wire[15:0] addr_remain3_750;
address_decode_4 decoder_3_750 = address_decode_4(addr_selector2_46[14],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_750,addr_remain3_750);


wire[15:0] addr_selector3_751;
wire[15:0] addr_remain3_751;
address_decode_4 decoder_3_751 = address_decode_4(addr_selector2_46[15],addr_remain2_46[15:0],addr_remain2_46,addr_selector3_751,addr_remain3_751);


wire[15:0] addr_selector3_752;
wire[15:0] addr_remain3_752;
address_decode_4 decoder_3_752 = address_decode_4(addr_selector2_47[0],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_752,addr_remain3_752);


wire[15:0] addr_selector3_753;
wire[15:0] addr_remain3_753;
address_decode_4 decoder_3_753 = address_decode_4(addr_selector2_47[1],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_753,addr_remain3_753);


wire[15:0] addr_selector3_754;
wire[15:0] addr_remain3_754;
address_decode_4 decoder_3_754 = address_decode_4(addr_selector2_47[2],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_754,addr_remain3_754);


wire[15:0] addr_selector3_755;
wire[15:0] addr_remain3_755;
address_decode_4 decoder_3_755 = address_decode_4(addr_selector2_47[3],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_755,addr_remain3_755);


wire[15:0] addr_selector3_756;
wire[15:0] addr_remain3_756;
address_decode_4 decoder_3_756 = address_decode_4(addr_selector2_47[4],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_756,addr_remain3_756);


wire[15:0] addr_selector3_757;
wire[15:0] addr_remain3_757;
address_decode_4 decoder_3_757 = address_decode_4(addr_selector2_47[5],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_757,addr_remain3_757);


wire[15:0] addr_selector3_758;
wire[15:0] addr_remain3_758;
address_decode_4 decoder_3_758 = address_decode_4(addr_selector2_47[6],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_758,addr_remain3_758);


wire[15:0] addr_selector3_759;
wire[15:0] addr_remain3_759;
address_decode_4 decoder_3_759 = address_decode_4(addr_selector2_47[7],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_759,addr_remain3_759);


wire[15:0] addr_selector3_760;
wire[15:0] addr_remain3_760;
address_decode_4 decoder_3_760 = address_decode_4(addr_selector2_47[8],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_760,addr_remain3_760);


wire[15:0] addr_selector3_761;
wire[15:0] addr_remain3_761;
address_decode_4 decoder_3_761 = address_decode_4(addr_selector2_47[9],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_761,addr_remain3_761);


wire[15:0] addr_selector3_762;
wire[15:0] addr_remain3_762;
address_decode_4 decoder_3_762 = address_decode_4(addr_selector2_47[10],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_762,addr_remain3_762);


wire[15:0] addr_selector3_763;
wire[15:0] addr_remain3_763;
address_decode_4 decoder_3_763 = address_decode_4(addr_selector2_47[11],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_763,addr_remain3_763);


wire[15:0] addr_selector3_764;
wire[15:0] addr_remain3_764;
address_decode_4 decoder_3_764 = address_decode_4(addr_selector2_47[12],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_764,addr_remain3_764);


wire[15:0] addr_selector3_765;
wire[15:0] addr_remain3_765;
address_decode_4 decoder_3_765 = address_decode_4(addr_selector2_47[13],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_765,addr_remain3_765);


wire[15:0] addr_selector3_766;
wire[15:0] addr_remain3_766;
address_decode_4 decoder_3_766 = address_decode_4(addr_selector2_47[14],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_766,addr_remain3_766);


wire[15:0] addr_selector3_767;
wire[15:0] addr_remain3_767;
address_decode_4 decoder_3_767 = address_decode_4(addr_selector2_47[15],addr_remain2_47[15:0],addr_remain2_47,addr_selector3_767,addr_remain3_767);


wire[15:0] addr_selector3_768;
wire[15:0] addr_remain3_768;
address_decode_4 decoder_3_768 = address_decode_4(addr_selector2_48[0],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_768,addr_remain3_768);


wire[15:0] addr_selector3_769;
wire[15:0] addr_remain3_769;
address_decode_4 decoder_3_769 = address_decode_4(addr_selector2_48[1],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_769,addr_remain3_769);


wire[15:0] addr_selector3_770;
wire[15:0] addr_remain3_770;
address_decode_4 decoder_3_770 = address_decode_4(addr_selector2_48[2],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_770,addr_remain3_770);


wire[15:0] addr_selector3_771;
wire[15:0] addr_remain3_771;
address_decode_4 decoder_3_771 = address_decode_4(addr_selector2_48[3],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_771,addr_remain3_771);


wire[15:0] addr_selector3_772;
wire[15:0] addr_remain3_772;
address_decode_4 decoder_3_772 = address_decode_4(addr_selector2_48[4],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_772,addr_remain3_772);


wire[15:0] addr_selector3_773;
wire[15:0] addr_remain3_773;
address_decode_4 decoder_3_773 = address_decode_4(addr_selector2_48[5],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_773,addr_remain3_773);


wire[15:0] addr_selector3_774;
wire[15:0] addr_remain3_774;
address_decode_4 decoder_3_774 = address_decode_4(addr_selector2_48[6],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_774,addr_remain3_774);


wire[15:0] addr_selector3_775;
wire[15:0] addr_remain3_775;
address_decode_4 decoder_3_775 = address_decode_4(addr_selector2_48[7],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_775,addr_remain3_775);


wire[15:0] addr_selector3_776;
wire[15:0] addr_remain3_776;
address_decode_4 decoder_3_776 = address_decode_4(addr_selector2_48[8],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_776,addr_remain3_776);


wire[15:0] addr_selector3_777;
wire[15:0] addr_remain3_777;
address_decode_4 decoder_3_777 = address_decode_4(addr_selector2_48[9],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_777,addr_remain3_777);


wire[15:0] addr_selector3_778;
wire[15:0] addr_remain3_778;
address_decode_4 decoder_3_778 = address_decode_4(addr_selector2_48[10],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_778,addr_remain3_778);


wire[15:0] addr_selector3_779;
wire[15:0] addr_remain3_779;
address_decode_4 decoder_3_779 = address_decode_4(addr_selector2_48[11],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_779,addr_remain3_779);


wire[15:0] addr_selector3_780;
wire[15:0] addr_remain3_780;
address_decode_4 decoder_3_780 = address_decode_4(addr_selector2_48[12],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_780,addr_remain3_780);


wire[15:0] addr_selector3_781;
wire[15:0] addr_remain3_781;
address_decode_4 decoder_3_781 = address_decode_4(addr_selector2_48[13],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_781,addr_remain3_781);


wire[15:0] addr_selector3_782;
wire[15:0] addr_remain3_782;
address_decode_4 decoder_3_782 = address_decode_4(addr_selector2_48[14],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_782,addr_remain3_782);


wire[15:0] addr_selector3_783;
wire[15:0] addr_remain3_783;
address_decode_4 decoder_3_783 = address_decode_4(addr_selector2_48[15],addr_remain2_48[15:0],addr_remain2_48,addr_selector3_783,addr_remain3_783);


wire[15:0] addr_selector3_784;
wire[15:0] addr_remain3_784;
address_decode_4 decoder_3_784 = address_decode_4(addr_selector2_49[0],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_784,addr_remain3_784);


wire[15:0] addr_selector3_785;
wire[15:0] addr_remain3_785;
address_decode_4 decoder_3_785 = address_decode_4(addr_selector2_49[1],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_785,addr_remain3_785);


wire[15:0] addr_selector3_786;
wire[15:0] addr_remain3_786;
address_decode_4 decoder_3_786 = address_decode_4(addr_selector2_49[2],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_786,addr_remain3_786);


wire[15:0] addr_selector3_787;
wire[15:0] addr_remain3_787;
address_decode_4 decoder_3_787 = address_decode_4(addr_selector2_49[3],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_787,addr_remain3_787);


wire[15:0] addr_selector3_788;
wire[15:0] addr_remain3_788;
address_decode_4 decoder_3_788 = address_decode_4(addr_selector2_49[4],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_788,addr_remain3_788);


wire[15:0] addr_selector3_789;
wire[15:0] addr_remain3_789;
address_decode_4 decoder_3_789 = address_decode_4(addr_selector2_49[5],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_789,addr_remain3_789);


wire[15:0] addr_selector3_790;
wire[15:0] addr_remain3_790;
address_decode_4 decoder_3_790 = address_decode_4(addr_selector2_49[6],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_790,addr_remain3_790);


wire[15:0] addr_selector3_791;
wire[15:0] addr_remain3_791;
address_decode_4 decoder_3_791 = address_decode_4(addr_selector2_49[7],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_791,addr_remain3_791);


wire[15:0] addr_selector3_792;
wire[15:0] addr_remain3_792;
address_decode_4 decoder_3_792 = address_decode_4(addr_selector2_49[8],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_792,addr_remain3_792);


wire[15:0] addr_selector3_793;
wire[15:0] addr_remain3_793;
address_decode_4 decoder_3_793 = address_decode_4(addr_selector2_49[9],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_793,addr_remain3_793);


wire[15:0] addr_selector3_794;
wire[15:0] addr_remain3_794;
address_decode_4 decoder_3_794 = address_decode_4(addr_selector2_49[10],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_794,addr_remain3_794);


wire[15:0] addr_selector3_795;
wire[15:0] addr_remain3_795;
address_decode_4 decoder_3_795 = address_decode_4(addr_selector2_49[11],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_795,addr_remain3_795);


wire[15:0] addr_selector3_796;
wire[15:0] addr_remain3_796;
address_decode_4 decoder_3_796 = address_decode_4(addr_selector2_49[12],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_796,addr_remain3_796);


wire[15:0] addr_selector3_797;
wire[15:0] addr_remain3_797;
address_decode_4 decoder_3_797 = address_decode_4(addr_selector2_49[13],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_797,addr_remain3_797);


wire[15:0] addr_selector3_798;
wire[15:0] addr_remain3_798;
address_decode_4 decoder_3_798 = address_decode_4(addr_selector2_49[14],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_798,addr_remain3_798);


wire[15:0] addr_selector3_799;
wire[15:0] addr_remain3_799;
address_decode_4 decoder_3_799 = address_decode_4(addr_selector2_49[15],addr_remain2_49[15:0],addr_remain2_49,addr_selector3_799,addr_remain3_799);


wire[15:0] addr_selector3_800;
wire[15:0] addr_remain3_800;
address_decode_4 decoder_3_800 = address_decode_4(addr_selector2_50[0],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_800,addr_remain3_800);


wire[15:0] addr_selector3_801;
wire[15:0] addr_remain3_801;
address_decode_4 decoder_3_801 = address_decode_4(addr_selector2_50[1],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_801,addr_remain3_801);


wire[15:0] addr_selector3_802;
wire[15:0] addr_remain3_802;
address_decode_4 decoder_3_802 = address_decode_4(addr_selector2_50[2],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_802,addr_remain3_802);


wire[15:0] addr_selector3_803;
wire[15:0] addr_remain3_803;
address_decode_4 decoder_3_803 = address_decode_4(addr_selector2_50[3],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_803,addr_remain3_803);


wire[15:0] addr_selector3_804;
wire[15:0] addr_remain3_804;
address_decode_4 decoder_3_804 = address_decode_4(addr_selector2_50[4],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_804,addr_remain3_804);


wire[15:0] addr_selector3_805;
wire[15:0] addr_remain3_805;
address_decode_4 decoder_3_805 = address_decode_4(addr_selector2_50[5],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_805,addr_remain3_805);


wire[15:0] addr_selector3_806;
wire[15:0] addr_remain3_806;
address_decode_4 decoder_3_806 = address_decode_4(addr_selector2_50[6],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_806,addr_remain3_806);


wire[15:0] addr_selector3_807;
wire[15:0] addr_remain3_807;
address_decode_4 decoder_3_807 = address_decode_4(addr_selector2_50[7],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_807,addr_remain3_807);


wire[15:0] addr_selector3_808;
wire[15:0] addr_remain3_808;
address_decode_4 decoder_3_808 = address_decode_4(addr_selector2_50[8],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_808,addr_remain3_808);


wire[15:0] addr_selector3_809;
wire[15:0] addr_remain3_809;
address_decode_4 decoder_3_809 = address_decode_4(addr_selector2_50[9],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_809,addr_remain3_809);


wire[15:0] addr_selector3_810;
wire[15:0] addr_remain3_810;
address_decode_4 decoder_3_810 = address_decode_4(addr_selector2_50[10],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_810,addr_remain3_810);


wire[15:0] addr_selector3_811;
wire[15:0] addr_remain3_811;
address_decode_4 decoder_3_811 = address_decode_4(addr_selector2_50[11],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_811,addr_remain3_811);


wire[15:0] addr_selector3_812;
wire[15:0] addr_remain3_812;
address_decode_4 decoder_3_812 = address_decode_4(addr_selector2_50[12],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_812,addr_remain3_812);


wire[15:0] addr_selector3_813;
wire[15:0] addr_remain3_813;
address_decode_4 decoder_3_813 = address_decode_4(addr_selector2_50[13],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_813,addr_remain3_813);


wire[15:0] addr_selector3_814;
wire[15:0] addr_remain3_814;
address_decode_4 decoder_3_814 = address_decode_4(addr_selector2_50[14],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_814,addr_remain3_814);


wire[15:0] addr_selector3_815;
wire[15:0] addr_remain3_815;
address_decode_4 decoder_3_815 = address_decode_4(addr_selector2_50[15],addr_remain2_50[15:0],addr_remain2_50,addr_selector3_815,addr_remain3_815);


wire[15:0] addr_selector3_816;
wire[15:0] addr_remain3_816;
address_decode_4 decoder_3_816 = address_decode_4(addr_selector2_51[0],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_816,addr_remain3_816);


wire[15:0] addr_selector3_817;
wire[15:0] addr_remain3_817;
address_decode_4 decoder_3_817 = address_decode_4(addr_selector2_51[1],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_817,addr_remain3_817);


wire[15:0] addr_selector3_818;
wire[15:0] addr_remain3_818;
address_decode_4 decoder_3_818 = address_decode_4(addr_selector2_51[2],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_818,addr_remain3_818);


wire[15:0] addr_selector3_819;
wire[15:0] addr_remain3_819;
address_decode_4 decoder_3_819 = address_decode_4(addr_selector2_51[3],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_819,addr_remain3_819);


wire[15:0] addr_selector3_820;
wire[15:0] addr_remain3_820;
address_decode_4 decoder_3_820 = address_decode_4(addr_selector2_51[4],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_820,addr_remain3_820);


wire[15:0] addr_selector3_821;
wire[15:0] addr_remain3_821;
address_decode_4 decoder_3_821 = address_decode_4(addr_selector2_51[5],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_821,addr_remain3_821);


wire[15:0] addr_selector3_822;
wire[15:0] addr_remain3_822;
address_decode_4 decoder_3_822 = address_decode_4(addr_selector2_51[6],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_822,addr_remain3_822);


wire[15:0] addr_selector3_823;
wire[15:0] addr_remain3_823;
address_decode_4 decoder_3_823 = address_decode_4(addr_selector2_51[7],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_823,addr_remain3_823);


wire[15:0] addr_selector3_824;
wire[15:0] addr_remain3_824;
address_decode_4 decoder_3_824 = address_decode_4(addr_selector2_51[8],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_824,addr_remain3_824);


wire[15:0] addr_selector3_825;
wire[15:0] addr_remain3_825;
address_decode_4 decoder_3_825 = address_decode_4(addr_selector2_51[9],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_825,addr_remain3_825);


wire[15:0] addr_selector3_826;
wire[15:0] addr_remain3_826;
address_decode_4 decoder_3_826 = address_decode_4(addr_selector2_51[10],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_826,addr_remain3_826);


wire[15:0] addr_selector3_827;
wire[15:0] addr_remain3_827;
address_decode_4 decoder_3_827 = address_decode_4(addr_selector2_51[11],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_827,addr_remain3_827);


wire[15:0] addr_selector3_828;
wire[15:0] addr_remain3_828;
address_decode_4 decoder_3_828 = address_decode_4(addr_selector2_51[12],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_828,addr_remain3_828);


wire[15:0] addr_selector3_829;
wire[15:0] addr_remain3_829;
address_decode_4 decoder_3_829 = address_decode_4(addr_selector2_51[13],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_829,addr_remain3_829);


wire[15:0] addr_selector3_830;
wire[15:0] addr_remain3_830;
address_decode_4 decoder_3_830 = address_decode_4(addr_selector2_51[14],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_830,addr_remain3_830);


wire[15:0] addr_selector3_831;
wire[15:0] addr_remain3_831;
address_decode_4 decoder_3_831 = address_decode_4(addr_selector2_51[15],addr_remain2_51[15:0],addr_remain2_51,addr_selector3_831,addr_remain3_831);


wire[15:0] addr_selector3_832;
wire[15:0] addr_remain3_832;
address_decode_4 decoder_3_832 = address_decode_4(addr_selector2_52[0],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_832,addr_remain3_832);


wire[15:0] addr_selector3_833;
wire[15:0] addr_remain3_833;
address_decode_4 decoder_3_833 = address_decode_4(addr_selector2_52[1],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_833,addr_remain3_833);


wire[15:0] addr_selector3_834;
wire[15:0] addr_remain3_834;
address_decode_4 decoder_3_834 = address_decode_4(addr_selector2_52[2],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_834,addr_remain3_834);


wire[15:0] addr_selector3_835;
wire[15:0] addr_remain3_835;
address_decode_4 decoder_3_835 = address_decode_4(addr_selector2_52[3],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_835,addr_remain3_835);


wire[15:0] addr_selector3_836;
wire[15:0] addr_remain3_836;
address_decode_4 decoder_3_836 = address_decode_4(addr_selector2_52[4],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_836,addr_remain3_836);


wire[15:0] addr_selector3_837;
wire[15:0] addr_remain3_837;
address_decode_4 decoder_3_837 = address_decode_4(addr_selector2_52[5],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_837,addr_remain3_837);


wire[15:0] addr_selector3_838;
wire[15:0] addr_remain3_838;
address_decode_4 decoder_3_838 = address_decode_4(addr_selector2_52[6],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_838,addr_remain3_838);


wire[15:0] addr_selector3_839;
wire[15:0] addr_remain3_839;
address_decode_4 decoder_3_839 = address_decode_4(addr_selector2_52[7],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_839,addr_remain3_839);


wire[15:0] addr_selector3_840;
wire[15:0] addr_remain3_840;
address_decode_4 decoder_3_840 = address_decode_4(addr_selector2_52[8],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_840,addr_remain3_840);


wire[15:0] addr_selector3_841;
wire[15:0] addr_remain3_841;
address_decode_4 decoder_3_841 = address_decode_4(addr_selector2_52[9],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_841,addr_remain3_841);


wire[15:0] addr_selector3_842;
wire[15:0] addr_remain3_842;
address_decode_4 decoder_3_842 = address_decode_4(addr_selector2_52[10],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_842,addr_remain3_842);


wire[15:0] addr_selector3_843;
wire[15:0] addr_remain3_843;
address_decode_4 decoder_3_843 = address_decode_4(addr_selector2_52[11],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_843,addr_remain3_843);


wire[15:0] addr_selector3_844;
wire[15:0] addr_remain3_844;
address_decode_4 decoder_3_844 = address_decode_4(addr_selector2_52[12],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_844,addr_remain3_844);


wire[15:0] addr_selector3_845;
wire[15:0] addr_remain3_845;
address_decode_4 decoder_3_845 = address_decode_4(addr_selector2_52[13],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_845,addr_remain3_845);


wire[15:0] addr_selector3_846;
wire[15:0] addr_remain3_846;
address_decode_4 decoder_3_846 = address_decode_4(addr_selector2_52[14],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_846,addr_remain3_846);


wire[15:0] addr_selector3_847;
wire[15:0] addr_remain3_847;
address_decode_4 decoder_3_847 = address_decode_4(addr_selector2_52[15],addr_remain2_52[15:0],addr_remain2_52,addr_selector3_847,addr_remain3_847);


wire[15:0] addr_selector3_848;
wire[15:0] addr_remain3_848;
address_decode_4 decoder_3_848 = address_decode_4(addr_selector2_53[0],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_848,addr_remain3_848);


wire[15:0] addr_selector3_849;
wire[15:0] addr_remain3_849;
address_decode_4 decoder_3_849 = address_decode_4(addr_selector2_53[1],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_849,addr_remain3_849);


wire[15:0] addr_selector3_850;
wire[15:0] addr_remain3_850;
address_decode_4 decoder_3_850 = address_decode_4(addr_selector2_53[2],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_850,addr_remain3_850);


wire[15:0] addr_selector3_851;
wire[15:0] addr_remain3_851;
address_decode_4 decoder_3_851 = address_decode_4(addr_selector2_53[3],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_851,addr_remain3_851);


wire[15:0] addr_selector3_852;
wire[15:0] addr_remain3_852;
address_decode_4 decoder_3_852 = address_decode_4(addr_selector2_53[4],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_852,addr_remain3_852);


wire[15:0] addr_selector3_853;
wire[15:0] addr_remain3_853;
address_decode_4 decoder_3_853 = address_decode_4(addr_selector2_53[5],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_853,addr_remain3_853);


wire[15:0] addr_selector3_854;
wire[15:0] addr_remain3_854;
address_decode_4 decoder_3_854 = address_decode_4(addr_selector2_53[6],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_854,addr_remain3_854);


wire[15:0] addr_selector3_855;
wire[15:0] addr_remain3_855;
address_decode_4 decoder_3_855 = address_decode_4(addr_selector2_53[7],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_855,addr_remain3_855);


wire[15:0] addr_selector3_856;
wire[15:0] addr_remain3_856;
address_decode_4 decoder_3_856 = address_decode_4(addr_selector2_53[8],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_856,addr_remain3_856);


wire[15:0] addr_selector3_857;
wire[15:0] addr_remain3_857;
address_decode_4 decoder_3_857 = address_decode_4(addr_selector2_53[9],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_857,addr_remain3_857);


wire[15:0] addr_selector3_858;
wire[15:0] addr_remain3_858;
address_decode_4 decoder_3_858 = address_decode_4(addr_selector2_53[10],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_858,addr_remain3_858);


wire[15:0] addr_selector3_859;
wire[15:0] addr_remain3_859;
address_decode_4 decoder_3_859 = address_decode_4(addr_selector2_53[11],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_859,addr_remain3_859);


wire[15:0] addr_selector3_860;
wire[15:0] addr_remain3_860;
address_decode_4 decoder_3_860 = address_decode_4(addr_selector2_53[12],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_860,addr_remain3_860);


wire[15:0] addr_selector3_861;
wire[15:0] addr_remain3_861;
address_decode_4 decoder_3_861 = address_decode_4(addr_selector2_53[13],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_861,addr_remain3_861);


wire[15:0] addr_selector3_862;
wire[15:0] addr_remain3_862;
address_decode_4 decoder_3_862 = address_decode_4(addr_selector2_53[14],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_862,addr_remain3_862);


wire[15:0] addr_selector3_863;
wire[15:0] addr_remain3_863;
address_decode_4 decoder_3_863 = address_decode_4(addr_selector2_53[15],addr_remain2_53[15:0],addr_remain2_53,addr_selector3_863,addr_remain3_863);


wire[15:0] addr_selector3_864;
wire[15:0] addr_remain3_864;
address_decode_4 decoder_3_864 = address_decode_4(addr_selector2_54[0],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_864,addr_remain3_864);


wire[15:0] addr_selector3_865;
wire[15:0] addr_remain3_865;
address_decode_4 decoder_3_865 = address_decode_4(addr_selector2_54[1],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_865,addr_remain3_865);


wire[15:0] addr_selector3_866;
wire[15:0] addr_remain3_866;
address_decode_4 decoder_3_866 = address_decode_4(addr_selector2_54[2],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_866,addr_remain3_866);


wire[15:0] addr_selector3_867;
wire[15:0] addr_remain3_867;
address_decode_4 decoder_3_867 = address_decode_4(addr_selector2_54[3],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_867,addr_remain3_867);


wire[15:0] addr_selector3_868;
wire[15:0] addr_remain3_868;
address_decode_4 decoder_3_868 = address_decode_4(addr_selector2_54[4],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_868,addr_remain3_868);


wire[15:0] addr_selector3_869;
wire[15:0] addr_remain3_869;
address_decode_4 decoder_3_869 = address_decode_4(addr_selector2_54[5],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_869,addr_remain3_869);


wire[15:0] addr_selector3_870;
wire[15:0] addr_remain3_870;
address_decode_4 decoder_3_870 = address_decode_4(addr_selector2_54[6],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_870,addr_remain3_870);


wire[15:0] addr_selector3_871;
wire[15:0] addr_remain3_871;
address_decode_4 decoder_3_871 = address_decode_4(addr_selector2_54[7],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_871,addr_remain3_871);


wire[15:0] addr_selector3_872;
wire[15:0] addr_remain3_872;
address_decode_4 decoder_3_872 = address_decode_4(addr_selector2_54[8],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_872,addr_remain3_872);


wire[15:0] addr_selector3_873;
wire[15:0] addr_remain3_873;
address_decode_4 decoder_3_873 = address_decode_4(addr_selector2_54[9],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_873,addr_remain3_873);


wire[15:0] addr_selector3_874;
wire[15:0] addr_remain3_874;
address_decode_4 decoder_3_874 = address_decode_4(addr_selector2_54[10],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_874,addr_remain3_874);


wire[15:0] addr_selector3_875;
wire[15:0] addr_remain3_875;
address_decode_4 decoder_3_875 = address_decode_4(addr_selector2_54[11],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_875,addr_remain3_875);


wire[15:0] addr_selector3_876;
wire[15:0] addr_remain3_876;
address_decode_4 decoder_3_876 = address_decode_4(addr_selector2_54[12],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_876,addr_remain3_876);


wire[15:0] addr_selector3_877;
wire[15:0] addr_remain3_877;
address_decode_4 decoder_3_877 = address_decode_4(addr_selector2_54[13],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_877,addr_remain3_877);


wire[15:0] addr_selector3_878;
wire[15:0] addr_remain3_878;
address_decode_4 decoder_3_878 = address_decode_4(addr_selector2_54[14],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_878,addr_remain3_878);


wire[15:0] addr_selector3_879;
wire[15:0] addr_remain3_879;
address_decode_4 decoder_3_879 = address_decode_4(addr_selector2_54[15],addr_remain2_54[15:0],addr_remain2_54,addr_selector3_879,addr_remain3_879);


wire[15:0] addr_selector3_880;
wire[15:0] addr_remain3_880;
address_decode_4 decoder_3_880 = address_decode_4(addr_selector2_55[0],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_880,addr_remain3_880);


wire[15:0] addr_selector3_881;
wire[15:0] addr_remain3_881;
address_decode_4 decoder_3_881 = address_decode_4(addr_selector2_55[1],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_881,addr_remain3_881);


wire[15:0] addr_selector3_882;
wire[15:0] addr_remain3_882;
address_decode_4 decoder_3_882 = address_decode_4(addr_selector2_55[2],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_882,addr_remain3_882);


wire[15:0] addr_selector3_883;
wire[15:0] addr_remain3_883;
address_decode_4 decoder_3_883 = address_decode_4(addr_selector2_55[3],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_883,addr_remain3_883);


wire[15:0] addr_selector3_884;
wire[15:0] addr_remain3_884;
address_decode_4 decoder_3_884 = address_decode_4(addr_selector2_55[4],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_884,addr_remain3_884);


wire[15:0] addr_selector3_885;
wire[15:0] addr_remain3_885;
address_decode_4 decoder_3_885 = address_decode_4(addr_selector2_55[5],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_885,addr_remain3_885);


wire[15:0] addr_selector3_886;
wire[15:0] addr_remain3_886;
address_decode_4 decoder_3_886 = address_decode_4(addr_selector2_55[6],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_886,addr_remain3_886);


wire[15:0] addr_selector3_887;
wire[15:0] addr_remain3_887;
address_decode_4 decoder_3_887 = address_decode_4(addr_selector2_55[7],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_887,addr_remain3_887);


wire[15:0] addr_selector3_888;
wire[15:0] addr_remain3_888;
address_decode_4 decoder_3_888 = address_decode_4(addr_selector2_55[8],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_888,addr_remain3_888);


wire[15:0] addr_selector3_889;
wire[15:0] addr_remain3_889;
address_decode_4 decoder_3_889 = address_decode_4(addr_selector2_55[9],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_889,addr_remain3_889);


wire[15:0] addr_selector3_890;
wire[15:0] addr_remain3_890;
address_decode_4 decoder_3_890 = address_decode_4(addr_selector2_55[10],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_890,addr_remain3_890);


wire[15:0] addr_selector3_891;
wire[15:0] addr_remain3_891;
address_decode_4 decoder_3_891 = address_decode_4(addr_selector2_55[11],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_891,addr_remain3_891);


wire[15:0] addr_selector3_892;
wire[15:0] addr_remain3_892;
address_decode_4 decoder_3_892 = address_decode_4(addr_selector2_55[12],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_892,addr_remain3_892);


wire[15:0] addr_selector3_893;
wire[15:0] addr_remain3_893;
address_decode_4 decoder_3_893 = address_decode_4(addr_selector2_55[13],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_893,addr_remain3_893);


wire[15:0] addr_selector3_894;
wire[15:0] addr_remain3_894;
address_decode_4 decoder_3_894 = address_decode_4(addr_selector2_55[14],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_894,addr_remain3_894);


wire[15:0] addr_selector3_895;
wire[15:0] addr_remain3_895;
address_decode_4 decoder_3_895 = address_decode_4(addr_selector2_55[15],addr_remain2_55[15:0],addr_remain2_55,addr_selector3_895,addr_remain3_895);


wire[15:0] addr_selector3_896;
wire[15:0] addr_remain3_896;
address_decode_4 decoder_3_896 = address_decode_4(addr_selector2_56[0],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_896,addr_remain3_896);


wire[15:0] addr_selector3_897;
wire[15:0] addr_remain3_897;
address_decode_4 decoder_3_897 = address_decode_4(addr_selector2_56[1],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_897,addr_remain3_897);


wire[15:0] addr_selector3_898;
wire[15:0] addr_remain3_898;
address_decode_4 decoder_3_898 = address_decode_4(addr_selector2_56[2],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_898,addr_remain3_898);


wire[15:0] addr_selector3_899;
wire[15:0] addr_remain3_899;
address_decode_4 decoder_3_899 = address_decode_4(addr_selector2_56[3],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_899,addr_remain3_899);


wire[15:0] addr_selector3_900;
wire[15:0] addr_remain3_900;
address_decode_4 decoder_3_900 = address_decode_4(addr_selector2_56[4],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_900,addr_remain3_900);


wire[15:0] addr_selector3_901;
wire[15:0] addr_remain3_901;
address_decode_4 decoder_3_901 = address_decode_4(addr_selector2_56[5],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_901,addr_remain3_901);


wire[15:0] addr_selector3_902;
wire[15:0] addr_remain3_902;
address_decode_4 decoder_3_902 = address_decode_4(addr_selector2_56[6],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_902,addr_remain3_902);


wire[15:0] addr_selector3_903;
wire[15:0] addr_remain3_903;
address_decode_4 decoder_3_903 = address_decode_4(addr_selector2_56[7],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_903,addr_remain3_903);


wire[15:0] addr_selector3_904;
wire[15:0] addr_remain3_904;
address_decode_4 decoder_3_904 = address_decode_4(addr_selector2_56[8],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_904,addr_remain3_904);


wire[15:0] addr_selector3_905;
wire[15:0] addr_remain3_905;
address_decode_4 decoder_3_905 = address_decode_4(addr_selector2_56[9],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_905,addr_remain3_905);


wire[15:0] addr_selector3_906;
wire[15:0] addr_remain3_906;
address_decode_4 decoder_3_906 = address_decode_4(addr_selector2_56[10],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_906,addr_remain3_906);


wire[15:0] addr_selector3_907;
wire[15:0] addr_remain3_907;
address_decode_4 decoder_3_907 = address_decode_4(addr_selector2_56[11],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_907,addr_remain3_907);


wire[15:0] addr_selector3_908;
wire[15:0] addr_remain3_908;
address_decode_4 decoder_3_908 = address_decode_4(addr_selector2_56[12],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_908,addr_remain3_908);


wire[15:0] addr_selector3_909;
wire[15:0] addr_remain3_909;
address_decode_4 decoder_3_909 = address_decode_4(addr_selector2_56[13],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_909,addr_remain3_909);


wire[15:0] addr_selector3_910;
wire[15:0] addr_remain3_910;
address_decode_4 decoder_3_910 = address_decode_4(addr_selector2_56[14],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_910,addr_remain3_910);


wire[15:0] addr_selector3_911;
wire[15:0] addr_remain3_911;
address_decode_4 decoder_3_911 = address_decode_4(addr_selector2_56[15],addr_remain2_56[15:0],addr_remain2_56,addr_selector3_911,addr_remain3_911);


wire[15:0] addr_selector3_912;
wire[15:0] addr_remain3_912;
address_decode_4 decoder_3_912 = address_decode_4(addr_selector2_57[0],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_912,addr_remain3_912);


wire[15:0] addr_selector3_913;
wire[15:0] addr_remain3_913;
address_decode_4 decoder_3_913 = address_decode_4(addr_selector2_57[1],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_913,addr_remain3_913);


wire[15:0] addr_selector3_914;
wire[15:0] addr_remain3_914;
address_decode_4 decoder_3_914 = address_decode_4(addr_selector2_57[2],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_914,addr_remain3_914);


wire[15:0] addr_selector3_915;
wire[15:0] addr_remain3_915;
address_decode_4 decoder_3_915 = address_decode_4(addr_selector2_57[3],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_915,addr_remain3_915);


wire[15:0] addr_selector3_916;
wire[15:0] addr_remain3_916;
address_decode_4 decoder_3_916 = address_decode_4(addr_selector2_57[4],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_916,addr_remain3_916);


wire[15:0] addr_selector3_917;
wire[15:0] addr_remain3_917;
address_decode_4 decoder_3_917 = address_decode_4(addr_selector2_57[5],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_917,addr_remain3_917);


wire[15:0] addr_selector3_918;
wire[15:0] addr_remain3_918;
address_decode_4 decoder_3_918 = address_decode_4(addr_selector2_57[6],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_918,addr_remain3_918);


wire[15:0] addr_selector3_919;
wire[15:0] addr_remain3_919;
address_decode_4 decoder_3_919 = address_decode_4(addr_selector2_57[7],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_919,addr_remain3_919);


wire[15:0] addr_selector3_920;
wire[15:0] addr_remain3_920;
address_decode_4 decoder_3_920 = address_decode_4(addr_selector2_57[8],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_920,addr_remain3_920);


wire[15:0] addr_selector3_921;
wire[15:0] addr_remain3_921;
address_decode_4 decoder_3_921 = address_decode_4(addr_selector2_57[9],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_921,addr_remain3_921);


wire[15:0] addr_selector3_922;
wire[15:0] addr_remain3_922;
address_decode_4 decoder_3_922 = address_decode_4(addr_selector2_57[10],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_922,addr_remain3_922);


wire[15:0] addr_selector3_923;
wire[15:0] addr_remain3_923;
address_decode_4 decoder_3_923 = address_decode_4(addr_selector2_57[11],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_923,addr_remain3_923);


wire[15:0] addr_selector3_924;
wire[15:0] addr_remain3_924;
address_decode_4 decoder_3_924 = address_decode_4(addr_selector2_57[12],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_924,addr_remain3_924);


wire[15:0] addr_selector3_925;
wire[15:0] addr_remain3_925;
address_decode_4 decoder_3_925 = address_decode_4(addr_selector2_57[13],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_925,addr_remain3_925);


wire[15:0] addr_selector3_926;
wire[15:0] addr_remain3_926;
address_decode_4 decoder_3_926 = address_decode_4(addr_selector2_57[14],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_926,addr_remain3_926);


wire[15:0] addr_selector3_927;
wire[15:0] addr_remain3_927;
address_decode_4 decoder_3_927 = address_decode_4(addr_selector2_57[15],addr_remain2_57[15:0],addr_remain2_57,addr_selector3_927,addr_remain3_927);


wire[15:0] addr_selector3_928;
wire[15:0] addr_remain3_928;
address_decode_4 decoder_3_928 = address_decode_4(addr_selector2_58[0],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_928,addr_remain3_928);


wire[15:0] addr_selector3_929;
wire[15:0] addr_remain3_929;
address_decode_4 decoder_3_929 = address_decode_4(addr_selector2_58[1],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_929,addr_remain3_929);


wire[15:0] addr_selector3_930;
wire[15:0] addr_remain3_930;
address_decode_4 decoder_3_930 = address_decode_4(addr_selector2_58[2],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_930,addr_remain3_930);


wire[15:0] addr_selector3_931;
wire[15:0] addr_remain3_931;
address_decode_4 decoder_3_931 = address_decode_4(addr_selector2_58[3],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_931,addr_remain3_931);


wire[15:0] addr_selector3_932;
wire[15:0] addr_remain3_932;
address_decode_4 decoder_3_932 = address_decode_4(addr_selector2_58[4],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_932,addr_remain3_932);


wire[15:0] addr_selector3_933;
wire[15:0] addr_remain3_933;
address_decode_4 decoder_3_933 = address_decode_4(addr_selector2_58[5],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_933,addr_remain3_933);


wire[15:0] addr_selector3_934;
wire[15:0] addr_remain3_934;
address_decode_4 decoder_3_934 = address_decode_4(addr_selector2_58[6],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_934,addr_remain3_934);


wire[15:0] addr_selector3_935;
wire[15:0] addr_remain3_935;
address_decode_4 decoder_3_935 = address_decode_4(addr_selector2_58[7],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_935,addr_remain3_935);


wire[15:0] addr_selector3_936;
wire[15:0] addr_remain3_936;
address_decode_4 decoder_3_936 = address_decode_4(addr_selector2_58[8],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_936,addr_remain3_936);


wire[15:0] addr_selector3_937;
wire[15:0] addr_remain3_937;
address_decode_4 decoder_3_937 = address_decode_4(addr_selector2_58[9],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_937,addr_remain3_937);


wire[15:0] addr_selector3_938;
wire[15:0] addr_remain3_938;
address_decode_4 decoder_3_938 = address_decode_4(addr_selector2_58[10],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_938,addr_remain3_938);


wire[15:0] addr_selector3_939;
wire[15:0] addr_remain3_939;
address_decode_4 decoder_3_939 = address_decode_4(addr_selector2_58[11],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_939,addr_remain3_939);


wire[15:0] addr_selector3_940;
wire[15:0] addr_remain3_940;
address_decode_4 decoder_3_940 = address_decode_4(addr_selector2_58[12],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_940,addr_remain3_940);


wire[15:0] addr_selector3_941;
wire[15:0] addr_remain3_941;
address_decode_4 decoder_3_941 = address_decode_4(addr_selector2_58[13],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_941,addr_remain3_941);


wire[15:0] addr_selector3_942;
wire[15:0] addr_remain3_942;
address_decode_4 decoder_3_942 = address_decode_4(addr_selector2_58[14],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_942,addr_remain3_942);


wire[15:0] addr_selector3_943;
wire[15:0] addr_remain3_943;
address_decode_4 decoder_3_943 = address_decode_4(addr_selector2_58[15],addr_remain2_58[15:0],addr_remain2_58,addr_selector3_943,addr_remain3_943);


wire[15:0] addr_selector3_944;
wire[15:0] addr_remain3_944;
address_decode_4 decoder_3_944 = address_decode_4(addr_selector2_59[0],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_944,addr_remain3_944);


wire[15:0] addr_selector3_945;
wire[15:0] addr_remain3_945;
address_decode_4 decoder_3_945 = address_decode_4(addr_selector2_59[1],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_945,addr_remain3_945);


wire[15:0] addr_selector3_946;
wire[15:0] addr_remain3_946;
address_decode_4 decoder_3_946 = address_decode_4(addr_selector2_59[2],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_946,addr_remain3_946);


wire[15:0] addr_selector3_947;
wire[15:0] addr_remain3_947;
address_decode_4 decoder_3_947 = address_decode_4(addr_selector2_59[3],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_947,addr_remain3_947);


wire[15:0] addr_selector3_948;
wire[15:0] addr_remain3_948;
address_decode_4 decoder_3_948 = address_decode_4(addr_selector2_59[4],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_948,addr_remain3_948);


wire[15:0] addr_selector3_949;
wire[15:0] addr_remain3_949;
address_decode_4 decoder_3_949 = address_decode_4(addr_selector2_59[5],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_949,addr_remain3_949);


wire[15:0] addr_selector3_950;
wire[15:0] addr_remain3_950;
address_decode_4 decoder_3_950 = address_decode_4(addr_selector2_59[6],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_950,addr_remain3_950);


wire[15:0] addr_selector3_951;
wire[15:0] addr_remain3_951;
address_decode_4 decoder_3_951 = address_decode_4(addr_selector2_59[7],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_951,addr_remain3_951);


wire[15:0] addr_selector3_952;
wire[15:0] addr_remain3_952;
address_decode_4 decoder_3_952 = address_decode_4(addr_selector2_59[8],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_952,addr_remain3_952);


wire[15:0] addr_selector3_953;
wire[15:0] addr_remain3_953;
address_decode_4 decoder_3_953 = address_decode_4(addr_selector2_59[9],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_953,addr_remain3_953);


wire[15:0] addr_selector3_954;
wire[15:0] addr_remain3_954;
address_decode_4 decoder_3_954 = address_decode_4(addr_selector2_59[10],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_954,addr_remain3_954);


wire[15:0] addr_selector3_955;
wire[15:0] addr_remain3_955;
address_decode_4 decoder_3_955 = address_decode_4(addr_selector2_59[11],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_955,addr_remain3_955);


wire[15:0] addr_selector3_956;
wire[15:0] addr_remain3_956;
address_decode_4 decoder_3_956 = address_decode_4(addr_selector2_59[12],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_956,addr_remain3_956);


wire[15:0] addr_selector3_957;
wire[15:0] addr_remain3_957;
address_decode_4 decoder_3_957 = address_decode_4(addr_selector2_59[13],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_957,addr_remain3_957);


wire[15:0] addr_selector3_958;
wire[15:0] addr_remain3_958;
address_decode_4 decoder_3_958 = address_decode_4(addr_selector2_59[14],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_958,addr_remain3_958);


wire[15:0] addr_selector3_959;
wire[15:0] addr_remain3_959;
address_decode_4 decoder_3_959 = address_decode_4(addr_selector2_59[15],addr_remain2_59[15:0],addr_remain2_59,addr_selector3_959,addr_remain3_959);


wire[15:0] addr_selector3_960;
wire[15:0] addr_remain3_960;
address_decode_4 decoder_3_960 = address_decode_4(addr_selector2_60[0],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_960,addr_remain3_960);


wire[15:0] addr_selector3_961;
wire[15:0] addr_remain3_961;
address_decode_4 decoder_3_961 = address_decode_4(addr_selector2_60[1],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_961,addr_remain3_961);


wire[15:0] addr_selector3_962;
wire[15:0] addr_remain3_962;
address_decode_4 decoder_3_962 = address_decode_4(addr_selector2_60[2],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_962,addr_remain3_962);


wire[15:0] addr_selector3_963;
wire[15:0] addr_remain3_963;
address_decode_4 decoder_3_963 = address_decode_4(addr_selector2_60[3],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_963,addr_remain3_963);


wire[15:0] addr_selector3_964;
wire[15:0] addr_remain3_964;
address_decode_4 decoder_3_964 = address_decode_4(addr_selector2_60[4],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_964,addr_remain3_964);


wire[15:0] addr_selector3_965;
wire[15:0] addr_remain3_965;
address_decode_4 decoder_3_965 = address_decode_4(addr_selector2_60[5],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_965,addr_remain3_965);


wire[15:0] addr_selector3_966;
wire[15:0] addr_remain3_966;
address_decode_4 decoder_3_966 = address_decode_4(addr_selector2_60[6],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_966,addr_remain3_966);


wire[15:0] addr_selector3_967;
wire[15:0] addr_remain3_967;
address_decode_4 decoder_3_967 = address_decode_4(addr_selector2_60[7],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_967,addr_remain3_967);


wire[15:0] addr_selector3_968;
wire[15:0] addr_remain3_968;
address_decode_4 decoder_3_968 = address_decode_4(addr_selector2_60[8],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_968,addr_remain3_968);


wire[15:0] addr_selector3_969;
wire[15:0] addr_remain3_969;
address_decode_4 decoder_3_969 = address_decode_4(addr_selector2_60[9],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_969,addr_remain3_969);


wire[15:0] addr_selector3_970;
wire[15:0] addr_remain3_970;
address_decode_4 decoder_3_970 = address_decode_4(addr_selector2_60[10],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_970,addr_remain3_970);


wire[15:0] addr_selector3_971;
wire[15:0] addr_remain3_971;
address_decode_4 decoder_3_971 = address_decode_4(addr_selector2_60[11],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_971,addr_remain3_971);


wire[15:0] addr_selector3_972;
wire[15:0] addr_remain3_972;
address_decode_4 decoder_3_972 = address_decode_4(addr_selector2_60[12],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_972,addr_remain3_972);


wire[15:0] addr_selector3_973;
wire[15:0] addr_remain3_973;
address_decode_4 decoder_3_973 = address_decode_4(addr_selector2_60[13],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_973,addr_remain3_973);


wire[15:0] addr_selector3_974;
wire[15:0] addr_remain3_974;
address_decode_4 decoder_3_974 = address_decode_4(addr_selector2_60[14],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_974,addr_remain3_974);


wire[15:0] addr_selector3_975;
wire[15:0] addr_remain3_975;
address_decode_4 decoder_3_975 = address_decode_4(addr_selector2_60[15],addr_remain2_60[15:0],addr_remain2_60,addr_selector3_975,addr_remain3_975);


wire[15:0] addr_selector3_976;
wire[15:0] addr_remain3_976;
address_decode_4 decoder_3_976 = address_decode_4(addr_selector2_61[0],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_976,addr_remain3_976);


wire[15:0] addr_selector3_977;
wire[15:0] addr_remain3_977;
address_decode_4 decoder_3_977 = address_decode_4(addr_selector2_61[1],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_977,addr_remain3_977);


wire[15:0] addr_selector3_978;
wire[15:0] addr_remain3_978;
address_decode_4 decoder_3_978 = address_decode_4(addr_selector2_61[2],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_978,addr_remain3_978);


wire[15:0] addr_selector3_979;
wire[15:0] addr_remain3_979;
address_decode_4 decoder_3_979 = address_decode_4(addr_selector2_61[3],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_979,addr_remain3_979);


wire[15:0] addr_selector3_980;
wire[15:0] addr_remain3_980;
address_decode_4 decoder_3_980 = address_decode_4(addr_selector2_61[4],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_980,addr_remain3_980);


wire[15:0] addr_selector3_981;
wire[15:0] addr_remain3_981;
address_decode_4 decoder_3_981 = address_decode_4(addr_selector2_61[5],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_981,addr_remain3_981);


wire[15:0] addr_selector3_982;
wire[15:0] addr_remain3_982;
address_decode_4 decoder_3_982 = address_decode_4(addr_selector2_61[6],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_982,addr_remain3_982);


wire[15:0] addr_selector3_983;
wire[15:0] addr_remain3_983;
address_decode_4 decoder_3_983 = address_decode_4(addr_selector2_61[7],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_983,addr_remain3_983);


wire[15:0] addr_selector3_984;
wire[15:0] addr_remain3_984;
address_decode_4 decoder_3_984 = address_decode_4(addr_selector2_61[8],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_984,addr_remain3_984);


wire[15:0] addr_selector3_985;
wire[15:0] addr_remain3_985;
address_decode_4 decoder_3_985 = address_decode_4(addr_selector2_61[9],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_985,addr_remain3_985);


wire[15:0] addr_selector3_986;
wire[15:0] addr_remain3_986;
address_decode_4 decoder_3_986 = address_decode_4(addr_selector2_61[10],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_986,addr_remain3_986);


wire[15:0] addr_selector3_987;
wire[15:0] addr_remain3_987;
address_decode_4 decoder_3_987 = address_decode_4(addr_selector2_61[11],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_987,addr_remain3_987);


wire[15:0] addr_selector3_988;
wire[15:0] addr_remain3_988;
address_decode_4 decoder_3_988 = address_decode_4(addr_selector2_61[12],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_988,addr_remain3_988);


wire[15:0] addr_selector3_989;
wire[15:0] addr_remain3_989;
address_decode_4 decoder_3_989 = address_decode_4(addr_selector2_61[13],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_989,addr_remain3_989);


wire[15:0] addr_selector3_990;
wire[15:0] addr_remain3_990;
address_decode_4 decoder_3_990 = address_decode_4(addr_selector2_61[14],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_990,addr_remain3_990);


wire[15:0] addr_selector3_991;
wire[15:0] addr_remain3_991;
address_decode_4 decoder_3_991 = address_decode_4(addr_selector2_61[15],addr_remain2_61[15:0],addr_remain2_61,addr_selector3_991,addr_remain3_991);


wire[15:0] addr_selector3_992;
wire[15:0] addr_remain3_992;
address_decode_4 decoder_3_992 = address_decode_4(addr_selector2_62[0],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_992,addr_remain3_992);


wire[15:0] addr_selector3_993;
wire[15:0] addr_remain3_993;
address_decode_4 decoder_3_993 = address_decode_4(addr_selector2_62[1],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_993,addr_remain3_993);


wire[15:0] addr_selector3_994;
wire[15:0] addr_remain3_994;
address_decode_4 decoder_3_994 = address_decode_4(addr_selector2_62[2],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_994,addr_remain3_994);


wire[15:0] addr_selector3_995;
wire[15:0] addr_remain3_995;
address_decode_4 decoder_3_995 = address_decode_4(addr_selector2_62[3],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_995,addr_remain3_995);


wire[15:0] addr_selector3_996;
wire[15:0] addr_remain3_996;
address_decode_4 decoder_3_996 = address_decode_4(addr_selector2_62[4],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_996,addr_remain3_996);


wire[15:0] addr_selector3_997;
wire[15:0] addr_remain3_997;
address_decode_4 decoder_3_997 = address_decode_4(addr_selector2_62[5],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_997,addr_remain3_997);


wire[15:0] addr_selector3_998;
wire[15:0] addr_remain3_998;
address_decode_4 decoder_3_998 = address_decode_4(addr_selector2_62[6],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_998,addr_remain3_998);


wire[15:0] addr_selector3_999;
wire[15:0] addr_remain3_999;
address_decode_4 decoder_3_999 = address_decode_4(addr_selector2_62[7],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_999,addr_remain3_999);


wire[15:0] addr_selector3_1000;
wire[15:0] addr_remain3_1000;
address_decode_4 decoder_3_1000 = address_decode_4(addr_selector2_62[8],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1000,addr_remain3_1000);


wire[15:0] addr_selector3_1001;
wire[15:0] addr_remain3_1001;
address_decode_4 decoder_3_1001 = address_decode_4(addr_selector2_62[9],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1001,addr_remain3_1001);


wire[15:0] addr_selector3_1002;
wire[15:0] addr_remain3_1002;
address_decode_4 decoder_3_1002 = address_decode_4(addr_selector2_62[10],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1002,addr_remain3_1002);


wire[15:0] addr_selector3_1003;
wire[15:0] addr_remain3_1003;
address_decode_4 decoder_3_1003 = address_decode_4(addr_selector2_62[11],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1003,addr_remain3_1003);


wire[15:0] addr_selector3_1004;
wire[15:0] addr_remain3_1004;
address_decode_4 decoder_3_1004 = address_decode_4(addr_selector2_62[12],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1004,addr_remain3_1004);


wire[15:0] addr_selector3_1005;
wire[15:0] addr_remain3_1005;
address_decode_4 decoder_3_1005 = address_decode_4(addr_selector2_62[13],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1005,addr_remain3_1005);


wire[15:0] addr_selector3_1006;
wire[15:0] addr_remain3_1006;
address_decode_4 decoder_3_1006 = address_decode_4(addr_selector2_62[14],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1006,addr_remain3_1006);


wire[15:0] addr_selector3_1007;
wire[15:0] addr_remain3_1007;
address_decode_4 decoder_3_1007 = address_decode_4(addr_selector2_62[15],addr_remain2_62[15:0],addr_remain2_62,addr_selector3_1007,addr_remain3_1007);


wire[15:0] addr_selector3_1008;
wire[15:0] addr_remain3_1008;
address_decode_4 decoder_3_1008 = address_decode_4(addr_selector2_63[0],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1008,addr_remain3_1008);


wire[15:0] addr_selector3_1009;
wire[15:0] addr_remain3_1009;
address_decode_4 decoder_3_1009 = address_decode_4(addr_selector2_63[1],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1009,addr_remain3_1009);


wire[15:0] addr_selector3_1010;
wire[15:0] addr_remain3_1010;
address_decode_4 decoder_3_1010 = address_decode_4(addr_selector2_63[2],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1010,addr_remain3_1010);


wire[15:0] addr_selector3_1011;
wire[15:0] addr_remain3_1011;
address_decode_4 decoder_3_1011 = address_decode_4(addr_selector2_63[3],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1011,addr_remain3_1011);


wire[15:0] addr_selector3_1012;
wire[15:0] addr_remain3_1012;
address_decode_4 decoder_3_1012 = address_decode_4(addr_selector2_63[4],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1012,addr_remain3_1012);


wire[15:0] addr_selector3_1013;
wire[15:0] addr_remain3_1013;
address_decode_4 decoder_3_1013 = address_decode_4(addr_selector2_63[5],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1013,addr_remain3_1013);


wire[15:0] addr_selector3_1014;
wire[15:0] addr_remain3_1014;
address_decode_4 decoder_3_1014 = address_decode_4(addr_selector2_63[6],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1014,addr_remain3_1014);


wire[15:0] addr_selector3_1015;
wire[15:0] addr_remain3_1015;
address_decode_4 decoder_3_1015 = address_decode_4(addr_selector2_63[7],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1015,addr_remain3_1015);


wire[15:0] addr_selector3_1016;
wire[15:0] addr_remain3_1016;
address_decode_4 decoder_3_1016 = address_decode_4(addr_selector2_63[8],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1016,addr_remain3_1016);


wire[15:0] addr_selector3_1017;
wire[15:0] addr_remain3_1017;
address_decode_4 decoder_3_1017 = address_decode_4(addr_selector2_63[9],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1017,addr_remain3_1017);


wire[15:0] addr_selector3_1018;
wire[15:0] addr_remain3_1018;
address_decode_4 decoder_3_1018 = address_decode_4(addr_selector2_63[10],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1018,addr_remain3_1018);


wire[15:0] addr_selector3_1019;
wire[15:0] addr_remain3_1019;
address_decode_4 decoder_3_1019 = address_decode_4(addr_selector2_63[11],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1019,addr_remain3_1019);


wire[15:0] addr_selector3_1020;
wire[15:0] addr_remain3_1020;
address_decode_4 decoder_3_1020 = address_decode_4(addr_selector2_63[12],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1020,addr_remain3_1020);


wire[15:0] addr_selector3_1021;
wire[15:0] addr_remain3_1021;
address_decode_4 decoder_3_1021 = address_decode_4(addr_selector2_63[13],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1021,addr_remain3_1021);


wire[15:0] addr_selector3_1022;
wire[15:0] addr_remain3_1022;
address_decode_4 decoder_3_1022 = address_decode_4(addr_selector2_63[14],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1022,addr_remain3_1022);


wire[15:0] addr_selector3_1023;
wire[15:0] addr_remain3_1023;
address_decode_4 decoder_3_1023 = address_decode_4(addr_selector2_63[15],addr_remain2_63[15:0],addr_remain2_63,addr_selector3_1023,addr_remain3_1023);


wire[15:0] addr_selector3_1024;
wire[15:0] addr_remain3_1024;
address_decode_4 decoder_3_1024 = address_decode_4(addr_selector2_64[0],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1024,addr_remain3_1024);


wire[15:0] addr_selector3_1025;
wire[15:0] addr_remain3_1025;
address_decode_4 decoder_3_1025 = address_decode_4(addr_selector2_64[1],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1025,addr_remain3_1025);


wire[15:0] addr_selector3_1026;
wire[15:0] addr_remain3_1026;
address_decode_4 decoder_3_1026 = address_decode_4(addr_selector2_64[2],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1026,addr_remain3_1026);


wire[15:0] addr_selector3_1027;
wire[15:0] addr_remain3_1027;
address_decode_4 decoder_3_1027 = address_decode_4(addr_selector2_64[3],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1027,addr_remain3_1027);


wire[15:0] addr_selector3_1028;
wire[15:0] addr_remain3_1028;
address_decode_4 decoder_3_1028 = address_decode_4(addr_selector2_64[4],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1028,addr_remain3_1028);


wire[15:0] addr_selector3_1029;
wire[15:0] addr_remain3_1029;
address_decode_4 decoder_3_1029 = address_decode_4(addr_selector2_64[5],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1029,addr_remain3_1029);


wire[15:0] addr_selector3_1030;
wire[15:0] addr_remain3_1030;
address_decode_4 decoder_3_1030 = address_decode_4(addr_selector2_64[6],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1030,addr_remain3_1030);


wire[15:0] addr_selector3_1031;
wire[15:0] addr_remain3_1031;
address_decode_4 decoder_3_1031 = address_decode_4(addr_selector2_64[7],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1031,addr_remain3_1031);


wire[15:0] addr_selector3_1032;
wire[15:0] addr_remain3_1032;
address_decode_4 decoder_3_1032 = address_decode_4(addr_selector2_64[8],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1032,addr_remain3_1032);


wire[15:0] addr_selector3_1033;
wire[15:0] addr_remain3_1033;
address_decode_4 decoder_3_1033 = address_decode_4(addr_selector2_64[9],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1033,addr_remain3_1033);


wire[15:0] addr_selector3_1034;
wire[15:0] addr_remain3_1034;
address_decode_4 decoder_3_1034 = address_decode_4(addr_selector2_64[10],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1034,addr_remain3_1034);


wire[15:0] addr_selector3_1035;
wire[15:0] addr_remain3_1035;
address_decode_4 decoder_3_1035 = address_decode_4(addr_selector2_64[11],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1035,addr_remain3_1035);


wire[15:0] addr_selector3_1036;
wire[15:0] addr_remain3_1036;
address_decode_4 decoder_3_1036 = address_decode_4(addr_selector2_64[12],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1036,addr_remain3_1036);


wire[15:0] addr_selector3_1037;
wire[15:0] addr_remain3_1037;
address_decode_4 decoder_3_1037 = address_decode_4(addr_selector2_64[13],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1037,addr_remain3_1037);


wire[15:0] addr_selector3_1038;
wire[15:0] addr_remain3_1038;
address_decode_4 decoder_3_1038 = address_decode_4(addr_selector2_64[14],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1038,addr_remain3_1038);


wire[15:0] addr_selector3_1039;
wire[15:0] addr_remain3_1039;
address_decode_4 decoder_3_1039 = address_decode_4(addr_selector2_64[15],addr_remain2_64[15:0],addr_remain2_64,addr_selector3_1039,addr_remain3_1039);


wire[15:0] addr_selector3_1040;
wire[15:0] addr_remain3_1040;
address_decode_4 decoder_3_1040 = address_decode_4(addr_selector2_65[0],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1040,addr_remain3_1040);


wire[15:0] addr_selector3_1041;
wire[15:0] addr_remain3_1041;
address_decode_4 decoder_3_1041 = address_decode_4(addr_selector2_65[1],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1041,addr_remain3_1041);


wire[15:0] addr_selector3_1042;
wire[15:0] addr_remain3_1042;
address_decode_4 decoder_3_1042 = address_decode_4(addr_selector2_65[2],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1042,addr_remain3_1042);


wire[15:0] addr_selector3_1043;
wire[15:0] addr_remain3_1043;
address_decode_4 decoder_3_1043 = address_decode_4(addr_selector2_65[3],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1043,addr_remain3_1043);


wire[15:0] addr_selector3_1044;
wire[15:0] addr_remain3_1044;
address_decode_4 decoder_3_1044 = address_decode_4(addr_selector2_65[4],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1044,addr_remain3_1044);


wire[15:0] addr_selector3_1045;
wire[15:0] addr_remain3_1045;
address_decode_4 decoder_3_1045 = address_decode_4(addr_selector2_65[5],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1045,addr_remain3_1045);


wire[15:0] addr_selector3_1046;
wire[15:0] addr_remain3_1046;
address_decode_4 decoder_3_1046 = address_decode_4(addr_selector2_65[6],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1046,addr_remain3_1046);


wire[15:0] addr_selector3_1047;
wire[15:0] addr_remain3_1047;
address_decode_4 decoder_3_1047 = address_decode_4(addr_selector2_65[7],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1047,addr_remain3_1047);


wire[15:0] addr_selector3_1048;
wire[15:0] addr_remain3_1048;
address_decode_4 decoder_3_1048 = address_decode_4(addr_selector2_65[8],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1048,addr_remain3_1048);


wire[15:0] addr_selector3_1049;
wire[15:0] addr_remain3_1049;
address_decode_4 decoder_3_1049 = address_decode_4(addr_selector2_65[9],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1049,addr_remain3_1049);


wire[15:0] addr_selector3_1050;
wire[15:0] addr_remain3_1050;
address_decode_4 decoder_3_1050 = address_decode_4(addr_selector2_65[10],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1050,addr_remain3_1050);


wire[15:0] addr_selector3_1051;
wire[15:0] addr_remain3_1051;
address_decode_4 decoder_3_1051 = address_decode_4(addr_selector2_65[11],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1051,addr_remain3_1051);


wire[15:0] addr_selector3_1052;
wire[15:0] addr_remain3_1052;
address_decode_4 decoder_3_1052 = address_decode_4(addr_selector2_65[12],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1052,addr_remain3_1052);


wire[15:0] addr_selector3_1053;
wire[15:0] addr_remain3_1053;
address_decode_4 decoder_3_1053 = address_decode_4(addr_selector2_65[13],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1053,addr_remain3_1053);


wire[15:0] addr_selector3_1054;
wire[15:0] addr_remain3_1054;
address_decode_4 decoder_3_1054 = address_decode_4(addr_selector2_65[14],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1054,addr_remain3_1054);


wire[15:0] addr_selector3_1055;
wire[15:0] addr_remain3_1055;
address_decode_4 decoder_3_1055 = address_decode_4(addr_selector2_65[15],addr_remain2_65[15:0],addr_remain2_65,addr_selector3_1055,addr_remain3_1055);


wire[15:0] addr_selector3_1056;
wire[15:0] addr_remain3_1056;
address_decode_4 decoder_3_1056 = address_decode_4(addr_selector2_66[0],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1056,addr_remain3_1056);


wire[15:0] addr_selector3_1057;
wire[15:0] addr_remain3_1057;
address_decode_4 decoder_3_1057 = address_decode_4(addr_selector2_66[1],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1057,addr_remain3_1057);


wire[15:0] addr_selector3_1058;
wire[15:0] addr_remain3_1058;
address_decode_4 decoder_3_1058 = address_decode_4(addr_selector2_66[2],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1058,addr_remain3_1058);


wire[15:0] addr_selector3_1059;
wire[15:0] addr_remain3_1059;
address_decode_4 decoder_3_1059 = address_decode_4(addr_selector2_66[3],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1059,addr_remain3_1059);


wire[15:0] addr_selector3_1060;
wire[15:0] addr_remain3_1060;
address_decode_4 decoder_3_1060 = address_decode_4(addr_selector2_66[4],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1060,addr_remain3_1060);


wire[15:0] addr_selector3_1061;
wire[15:0] addr_remain3_1061;
address_decode_4 decoder_3_1061 = address_decode_4(addr_selector2_66[5],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1061,addr_remain3_1061);


wire[15:0] addr_selector3_1062;
wire[15:0] addr_remain3_1062;
address_decode_4 decoder_3_1062 = address_decode_4(addr_selector2_66[6],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1062,addr_remain3_1062);


wire[15:0] addr_selector3_1063;
wire[15:0] addr_remain3_1063;
address_decode_4 decoder_3_1063 = address_decode_4(addr_selector2_66[7],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1063,addr_remain3_1063);


wire[15:0] addr_selector3_1064;
wire[15:0] addr_remain3_1064;
address_decode_4 decoder_3_1064 = address_decode_4(addr_selector2_66[8],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1064,addr_remain3_1064);


wire[15:0] addr_selector3_1065;
wire[15:0] addr_remain3_1065;
address_decode_4 decoder_3_1065 = address_decode_4(addr_selector2_66[9],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1065,addr_remain3_1065);


wire[15:0] addr_selector3_1066;
wire[15:0] addr_remain3_1066;
address_decode_4 decoder_3_1066 = address_decode_4(addr_selector2_66[10],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1066,addr_remain3_1066);


wire[15:0] addr_selector3_1067;
wire[15:0] addr_remain3_1067;
address_decode_4 decoder_3_1067 = address_decode_4(addr_selector2_66[11],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1067,addr_remain3_1067);


wire[15:0] addr_selector3_1068;
wire[15:0] addr_remain3_1068;
address_decode_4 decoder_3_1068 = address_decode_4(addr_selector2_66[12],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1068,addr_remain3_1068);


wire[15:0] addr_selector3_1069;
wire[15:0] addr_remain3_1069;
address_decode_4 decoder_3_1069 = address_decode_4(addr_selector2_66[13],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1069,addr_remain3_1069);


wire[15:0] addr_selector3_1070;
wire[15:0] addr_remain3_1070;
address_decode_4 decoder_3_1070 = address_decode_4(addr_selector2_66[14],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1070,addr_remain3_1070);


wire[15:0] addr_selector3_1071;
wire[15:0] addr_remain3_1071;
address_decode_4 decoder_3_1071 = address_decode_4(addr_selector2_66[15],addr_remain2_66[15:0],addr_remain2_66,addr_selector3_1071,addr_remain3_1071);


wire[15:0] addr_selector3_1072;
wire[15:0] addr_remain3_1072;
address_decode_4 decoder_3_1072 = address_decode_4(addr_selector2_67[0],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1072,addr_remain3_1072);


wire[15:0] addr_selector3_1073;
wire[15:0] addr_remain3_1073;
address_decode_4 decoder_3_1073 = address_decode_4(addr_selector2_67[1],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1073,addr_remain3_1073);


wire[15:0] addr_selector3_1074;
wire[15:0] addr_remain3_1074;
address_decode_4 decoder_3_1074 = address_decode_4(addr_selector2_67[2],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1074,addr_remain3_1074);


wire[15:0] addr_selector3_1075;
wire[15:0] addr_remain3_1075;
address_decode_4 decoder_3_1075 = address_decode_4(addr_selector2_67[3],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1075,addr_remain3_1075);


wire[15:0] addr_selector3_1076;
wire[15:0] addr_remain3_1076;
address_decode_4 decoder_3_1076 = address_decode_4(addr_selector2_67[4],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1076,addr_remain3_1076);


wire[15:0] addr_selector3_1077;
wire[15:0] addr_remain3_1077;
address_decode_4 decoder_3_1077 = address_decode_4(addr_selector2_67[5],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1077,addr_remain3_1077);


wire[15:0] addr_selector3_1078;
wire[15:0] addr_remain3_1078;
address_decode_4 decoder_3_1078 = address_decode_4(addr_selector2_67[6],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1078,addr_remain3_1078);


wire[15:0] addr_selector3_1079;
wire[15:0] addr_remain3_1079;
address_decode_4 decoder_3_1079 = address_decode_4(addr_selector2_67[7],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1079,addr_remain3_1079);


wire[15:0] addr_selector3_1080;
wire[15:0] addr_remain3_1080;
address_decode_4 decoder_3_1080 = address_decode_4(addr_selector2_67[8],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1080,addr_remain3_1080);


wire[15:0] addr_selector3_1081;
wire[15:0] addr_remain3_1081;
address_decode_4 decoder_3_1081 = address_decode_4(addr_selector2_67[9],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1081,addr_remain3_1081);


wire[15:0] addr_selector3_1082;
wire[15:0] addr_remain3_1082;
address_decode_4 decoder_3_1082 = address_decode_4(addr_selector2_67[10],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1082,addr_remain3_1082);


wire[15:0] addr_selector3_1083;
wire[15:0] addr_remain3_1083;
address_decode_4 decoder_3_1083 = address_decode_4(addr_selector2_67[11],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1083,addr_remain3_1083);


wire[15:0] addr_selector3_1084;
wire[15:0] addr_remain3_1084;
address_decode_4 decoder_3_1084 = address_decode_4(addr_selector2_67[12],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1084,addr_remain3_1084);


wire[15:0] addr_selector3_1085;
wire[15:0] addr_remain3_1085;
address_decode_4 decoder_3_1085 = address_decode_4(addr_selector2_67[13],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1085,addr_remain3_1085);


wire[15:0] addr_selector3_1086;
wire[15:0] addr_remain3_1086;
address_decode_4 decoder_3_1086 = address_decode_4(addr_selector2_67[14],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1086,addr_remain3_1086);


wire[15:0] addr_selector3_1087;
wire[15:0] addr_remain3_1087;
address_decode_4 decoder_3_1087 = address_decode_4(addr_selector2_67[15],addr_remain2_67[15:0],addr_remain2_67,addr_selector3_1087,addr_remain3_1087);


wire[15:0] addr_selector3_1088;
wire[15:0] addr_remain3_1088;
address_decode_4 decoder_3_1088 = address_decode_4(addr_selector2_68[0],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1088,addr_remain3_1088);


wire[15:0] addr_selector3_1089;
wire[15:0] addr_remain3_1089;
address_decode_4 decoder_3_1089 = address_decode_4(addr_selector2_68[1],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1089,addr_remain3_1089);


wire[15:0] addr_selector3_1090;
wire[15:0] addr_remain3_1090;
address_decode_4 decoder_3_1090 = address_decode_4(addr_selector2_68[2],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1090,addr_remain3_1090);


wire[15:0] addr_selector3_1091;
wire[15:0] addr_remain3_1091;
address_decode_4 decoder_3_1091 = address_decode_4(addr_selector2_68[3],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1091,addr_remain3_1091);


wire[15:0] addr_selector3_1092;
wire[15:0] addr_remain3_1092;
address_decode_4 decoder_3_1092 = address_decode_4(addr_selector2_68[4],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1092,addr_remain3_1092);


wire[15:0] addr_selector3_1093;
wire[15:0] addr_remain3_1093;
address_decode_4 decoder_3_1093 = address_decode_4(addr_selector2_68[5],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1093,addr_remain3_1093);


wire[15:0] addr_selector3_1094;
wire[15:0] addr_remain3_1094;
address_decode_4 decoder_3_1094 = address_decode_4(addr_selector2_68[6],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1094,addr_remain3_1094);


wire[15:0] addr_selector3_1095;
wire[15:0] addr_remain3_1095;
address_decode_4 decoder_3_1095 = address_decode_4(addr_selector2_68[7],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1095,addr_remain3_1095);


wire[15:0] addr_selector3_1096;
wire[15:0] addr_remain3_1096;
address_decode_4 decoder_3_1096 = address_decode_4(addr_selector2_68[8],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1096,addr_remain3_1096);


wire[15:0] addr_selector3_1097;
wire[15:0] addr_remain3_1097;
address_decode_4 decoder_3_1097 = address_decode_4(addr_selector2_68[9],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1097,addr_remain3_1097);


wire[15:0] addr_selector3_1098;
wire[15:0] addr_remain3_1098;
address_decode_4 decoder_3_1098 = address_decode_4(addr_selector2_68[10],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1098,addr_remain3_1098);


wire[15:0] addr_selector3_1099;
wire[15:0] addr_remain3_1099;
address_decode_4 decoder_3_1099 = address_decode_4(addr_selector2_68[11],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1099,addr_remain3_1099);


wire[15:0] addr_selector3_1100;
wire[15:0] addr_remain3_1100;
address_decode_4 decoder_3_1100 = address_decode_4(addr_selector2_68[12],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1100,addr_remain3_1100);


wire[15:0] addr_selector3_1101;
wire[15:0] addr_remain3_1101;
address_decode_4 decoder_3_1101 = address_decode_4(addr_selector2_68[13],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1101,addr_remain3_1101);


wire[15:0] addr_selector3_1102;
wire[15:0] addr_remain3_1102;
address_decode_4 decoder_3_1102 = address_decode_4(addr_selector2_68[14],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1102,addr_remain3_1102);


wire[15:0] addr_selector3_1103;
wire[15:0] addr_remain3_1103;
address_decode_4 decoder_3_1103 = address_decode_4(addr_selector2_68[15],addr_remain2_68[15:0],addr_remain2_68,addr_selector3_1103,addr_remain3_1103);


wire[15:0] addr_selector3_1104;
wire[15:0] addr_remain3_1104;
address_decode_4 decoder_3_1104 = address_decode_4(addr_selector2_69[0],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1104,addr_remain3_1104);


wire[15:0] addr_selector3_1105;
wire[15:0] addr_remain3_1105;
address_decode_4 decoder_3_1105 = address_decode_4(addr_selector2_69[1],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1105,addr_remain3_1105);


wire[15:0] addr_selector3_1106;
wire[15:0] addr_remain3_1106;
address_decode_4 decoder_3_1106 = address_decode_4(addr_selector2_69[2],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1106,addr_remain3_1106);


wire[15:0] addr_selector3_1107;
wire[15:0] addr_remain3_1107;
address_decode_4 decoder_3_1107 = address_decode_4(addr_selector2_69[3],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1107,addr_remain3_1107);


wire[15:0] addr_selector3_1108;
wire[15:0] addr_remain3_1108;
address_decode_4 decoder_3_1108 = address_decode_4(addr_selector2_69[4],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1108,addr_remain3_1108);


wire[15:0] addr_selector3_1109;
wire[15:0] addr_remain3_1109;
address_decode_4 decoder_3_1109 = address_decode_4(addr_selector2_69[5],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1109,addr_remain3_1109);


wire[15:0] addr_selector3_1110;
wire[15:0] addr_remain3_1110;
address_decode_4 decoder_3_1110 = address_decode_4(addr_selector2_69[6],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1110,addr_remain3_1110);


wire[15:0] addr_selector3_1111;
wire[15:0] addr_remain3_1111;
address_decode_4 decoder_3_1111 = address_decode_4(addr_selector2_69[7],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1111,addr_remain3_1111);


wire[15:0] addr_selector3_1112;
wire[15:0] addr_remain3_1112;
address_decode_4 decoder_3_1112 = address_decode_4(addr_selector2_69[8],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1112,addr_remain3_1112);


wire[15:0] addr_selector3_1113;
wire[15:0] addr_remain3_1113;
address_decode_4 decoder_3_1113 = address_decode_4(addr_selector2_69[9],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1113,addr_remain3_1113);


wire[15:0] addr_selector3_1114;
wire[15:0] addr_remain3_1114;
address_decode_4 decoder_3_1114 = address_decode_4(addr_selector2_69[10],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1114,addr_remain3_1114);


wire[15:0] addr_selector3_1115;
wire[15:0] addr_remain3_1115;
address_decode_4 decoder_3_1115 = address_decode_4(addr_selector2_69[11],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1115,addr_remain3_1115);


wire[15:0] addr_selector3_1116;
wire[15:0] addr_remain3_1116;
address_decode_4 decoder_3_1116 = address_decode_4(addr_selector2_69[12],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1116,addr_remain3_1116);


wire[15:0] addr_selector3_1117;
wire[15:0] addr_remain3_1117;
address_decode_4 decoder_3_1117 = address_decode_4(addr_selector2_69[13],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1117,addr_remain3_1117);


wire[15:0] addr_selector3_1118;
wire[15:0] addr_remain3_1118;
address_decode_4 decoder_3_1118 = address_decode_4(addr_selector2_69[14],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1118,addr_remain3_1118);


wire[15:0] addr_selector3_1119;
wire[15:0] addr_remain3_1119;
address_decode_4 decoder_3_1119 = address_decode_4(addr_selector2_69[15],addr_remain2_69[15:0],addr_remain2_69,addr_selector3_1119,addr_remain3_1119);


wire[15:0] addr_selector3_1120;
wire[15:0] addr_remain3_1120;
address_decode_4 decoder_3_1120 = address_decode_4(addr_selector2_70[0],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1120,addr_remain3_1120);


wire[15:0] addr_selector3_1121;
wire[15:0] addr_remain3_1121;
address_decode_4 decoder_3_1121 = address_decode_4(addr_selector2_70[1],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1121,addr_remain3_1121);


wire[15:0] addr_selector3_1122;
wire[15:0] addr_remain3_1122;
address_decode_4 decoder_3_1122 = address_decode_4(addr_selector2_70[2],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1122,addr_remain3_1122);


wire[15:0] addr_selector3_1123;
wire[15:0] addr_remain3_1123;
address_decode_4 decoder_3_1123 = address_decode_4(addr_selector2_70[3],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1123,addr_remain3_1123);


wire[15:0] addr_selector3_1124;
wire[15:0] addr_remain3_1124;
address_decode_4 decoder_3_1124 = address_decode_4(addr_selector2_70[4],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1124,addr_remain3_1124);


wire[15:0] addr_selector3_1125;
wire[15:0] addr_remain3_1125;
address_decode_4 decoder_3_1125 = address_decode_4(addr_selector2_70[5],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1125,addr_remain3_1125);


wire[15:0] addr_selector3_1126;
wire[15:0] addr_remain3_1126;
address_decode_4 decoder_3_1126 = address_decode_4(addr_selector2_70[6],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1126,addr_remain3_1126);


wire[15:0] addr_selector3_1127;
wire[15:0] addr_remain3_1127;
address_decode_4 decoder_3_1127 = address_decode_4(addr_selector2_70[7],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1127,addr_remain3_1127);


wire[15:0] addr_selector3_1128;
wire[15:0] addr_remain3_1128;
address_decode_4 decoder_3_1128 = address_decode_4(addr_selector2_70[8],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1128,addr_remain3_1128);


wire[15:0] addr_selector3_1129;
wire[15:0] addr_remain3_1129;
address_decode_4 decoder_3_1129 = address_decode_4(addr_selector2_70[9],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1129,addr_remain3_1129);


wire[15:0] addr_selector3_1130;
wire[15:0] addr_remain3_1130;
address_decode_4 decoder_3_1130 = address_decode_4(addr_selector2_70[10],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1130,addr_remain3_1130);


wire[15:0] addr_selector3_1131;
wire[15:0] addr_remain3_1131;
address_decode_4 decoder_3_1131 = address_decode_4(addr_selector2_70[11],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1131,addr_remain3_1131);


wire[15:0] addr_selector3_1132;
wire[15:0] addr_remain3_1132;
address_decode_4 decoder_3_1132 = address_decode_4(addr_selector2_70[12],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1132,addr_remain3_1132);


wire[15:0] addr_selector3_1133;
wire[15:0] addr_remain3_1133;
address_decode_4 decoder_3_1133 = address_decode_4(addr_selector2_70[13],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1133,addr_remain3_1133);


wire[15:0] addr_selector3_1134;
wire[15:0] addr_remain3_1134;
address_decode_4 decoder_3_1134 = address_decode_4(addr_selector2_70[14],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1134,addr_remain3_1134);


wire[15:0] addr_selector3_1135;
wire[15:0] addr_remain3_1135;
address_decode_4 decoder_3_1135 = address_decode_4(addr_selector2_70[15],addr_remain2_70[15:0],addr_remain2_70,addr_selector3_1135,addr_remain3_1135);


wire[15:0] addr_selector3_1136;
wire[15:0] addr_remain3_1136;
address_decode_4 decoder_3_1136 = address_decode_4(addr_selector2_71[0],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1136,addr_remain3_1136);


wire[15:0] addr_selector3_1137;
wire[15:0] addr_remain3_1137;
address_decode_4 decoder_3_1137 = address_decode_4(addr_selector2_71[1],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1137,addr_remain3_1137);


wire[15:0] addr_selector3_1138;
wire[15:0] addr_remain3_1138;
address_decode_4 decoder_3_1138 = address_decode_4(addr_selector2_71[2],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1138,addr_remain3_1138);


wire[15:0] addr_selector3_1139;
wire[15:0] addr_remain3_1139;
address_decode_4 decoder_3_1139 = address_decode_4(addr_selector2_71[3],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1139,addr_remain3_1139);


wire[15:0] addr_selector3_1140;
wire[15:0] addr_remain3_1140;
address_decode_4 decoder_3_1140 = address_decode_4(addr_selector2_71[4],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1140,addr_remain3_1140);


wire[15:0] addr_selector3_1141;
wire[15:0] addr_remain3_1141;
address_decode_4 decoder_3_1141 = address_decode_4(addr_selector2_71[5],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1141,addr_remain3_1141);


wire[15:0] addr_selector3_1142;
wire[15:0] addr_remain3_1142;
address_decode_4 decoder_3_1142 = address_decode_4(addr_selector2_71[6],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1142,addr_remain3_1142);


wire[15:0] addr_selector3_1143;
wire[15:0] addr_remain3_1143;
address_decode_4 decoder_3_1143 = address_decode_4(addr_selector2_71[7],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1143,addr_remain3_1143);


wire[15:0] addr_selector3_1144;
wire[15:0] addr_remain3_1144;
address_decode_4 decoder_3_1144 = address_decode_4(addr_selector2_71[8],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1144,addr_remain3_1144);


wire[15:0] addr_selector3_1145;
wire[15:0] addr_remain3_1145;
address_decode_4 decoder_3_1145 = address_decode_4(addr_selector2_71[9],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1145,addr_remain3_1145);


wire[15:0] addr_selector3_1146;
wire[15:0] addr_remain3_1146;
address_decode_4 decoder_3_1146 = address_decode_4(addr_selector2_71[10],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1146,addr_remain3_1146);


wire[15:0] addr_selector3_1147;
wire[15:0] addr_remain3_1147;
address_decode_4 decoder_3_1147 = address_decode_4(addr_selector2_71[11],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1147,addr_remain3_1147);


wire[15:0] addr_selector3_1148;
wire[15:0] addr_remain3_1148;
address_decode_4 decoder_3_1148 = address_decode_4(addr_selector2_71[12],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1148,addr_remain3_1148);


wire[15:0] addr_selector3_1149;
wire[15:0] addr_remain3_1149;
address_decode_4 decoder_3_1149 = address_decode_4(addr_selector2_71[13],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1149,addr_remain3_1149);


wire[15:0] addr_selector3_1150;
wire[15:0] addr_remain3_1150;
address_decode_4 decoder_3_1150 = address_decode_4(addr_selector2_71[14],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1150,addr_remain3_1150);


wire[15:0] addr_selector3_1151;
wire[15:0] addr_remain3_1151;
address_decode_4 decoder_3_1151 = address_decode_4(addr_selector2_71[15],addr_remain2_71[15:0],addr_remain2_71,addr_selector3_1151,addr_remain3_1151);


wire[15:0] addr_selector3_1152;
wire[15:0] addr_remain3_1152;
address_decode_4 decoder_3_1152 = address_decode_4(addr_selector2_72[0],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1152,addr_remain3_1152);


wire[15:0] addr_selector3_1153;
wire[15:0] addr_remain3_1153;
address_decode_4 decoder_3_1153 = address_decode_4(addr_selector2_72[1],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1153,addr_remain3_1153);


wire[15:0] addr_selector3_1154;
wire[15:0] addr_remain3_1154;
address_decode_4 decoder_3_1154 = address_decode_4(addr_selector2_72[2],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1154,addr_remain3_1154);


wire[15:0] addr_selector3_1155;
wire[15:0] addr_remain3_1155;
address_decode_4 decoder_3_1155 = address_decode_4(addr_selector2_72[3],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1155,addr_remain3_1155);


wire[15:0] addr_selector3_1156;
wire[15:0] addr_remain3_1156;
address_decode_4 decoder_3_1156 = address_decode_4(addr_selector2_72[4],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1156,addr_remain3_1156);


wire[15:0] addr_selector3_1157;
wire[15:0] addr_remain3_1157;
address_decode_4 decoder_3_1157 = address_decode_4(addr_selector2_72[5],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1157,addr_remain3_1157);


wire[15:0] addr_selector3_1158;
wire[15:0] addr_remain3_1158;
address_decode_4 decoder_3_1158 = address_decode_4(addr_selector2_72[6],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1158,addr_remain3_1158);


wire[15:0] addr_selector3_1159;
wire[15:0] addr_remain3_1159;
address_decode_4 decoder_3_1159 = address_decode_4(addr_selector2_72[7],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1159,addr_remain3_1159);


wire[15:0] addr_selector3_1160;
wire[15:0] addr_remain3_1160;
address_decode_4 decoder_3_1160 = address_decode_4(addr_selector2_72[8],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1160,addr_remain3_1160);


wire[15:0] addr_selector3_1161;
wire[15:0] addr_remain3_1161;
address_decode_4 decoder_3_1161 = address_decode_4(addr_selector2_72[9],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1161,addr_remain3_1161);


wire[15:0] addr_selector3_1162;
wire[15:0] addr_remain3_1162;
address_decode_4 decoder_3_1162 = address_decode_4(addr_selector2_72[10],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1162,addr_remain3_1162);


wire[15:0] addr_selector3_1163;
wire[15:0] addr_remain3_1163;
address_decode_4 decoder_3_1163 = address_decode_4(addr_selector2_72[11],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1163,addr_remain3_1163);


wire[15:0] addr_selector3_1164;
wire[15:0] addr_remain3_1164;
address_decode_4 decoder_3_1164 = address_decode_4(addr_selector2_72[12],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1164,addr_remain3_1164);


wire[15:0] addr_selector3_1165;
wire[15:0] addr_remain3_1165;
address_decode_4 decoder_3_1165 = address_decode_4(addr_selector2_72[13],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1165,addr_remain3_1165);


wire[15:0] addr_selector3_1166;
wire[15:0] addr_remain3_1166;
address_decode_4 decoder_3_1166 = address_decode_4(addr_selector2_72[14],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1166,addr_remain3_1166);


wire[15:0] addr_selector3_1167;
wire[15:0] addr_remain3_1167;
address_decode_4 decoder_3_1167 = address_decode_4(addr_selector2_72[15],addr_remain2_72[15:0],addr_remain2_72,addr_selector3_1167,addr_remain3_1167);


wire[15:0] addr_selector3_1168;
wire[15:0] addr_remain3_1168;
address_decode_4 decoder_3_1168 = address_decode_4(addr_selector2_73[0],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1168,addr_remain3_1168);


wire[15:0] addr_selector3_1169;
wire[15:0] addr_remain3_1169;
address_decode_4 decoder_3_1169 = address_decode_4(addr_selector2_73[1],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1169,addr_remain3_1169);


wire[15:0] addr_selector3_1170;
wire[15:0] addr_remain3_1170;
address_decode_4 decoder_3_1170 = address_decode_4(addr_selector2_73[2],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1170,addr_remain3_1170);


wire[15:0] addr_selector3_1171;
wire[15:0] addr_remain3_1171;
address_decode_4 decoder_3_1171 = address_decode_4(addr_selector2_73[3],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1171,addr_remain3_1171);


wire[15:0] addr_selector3_1172;
wire[15:0] addr_remain3_1172;
address_decode_4 decoder_3_1172 = address_decode_4(addr_selector2_73[4],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1172,addr_remain3_1172);


wire[15:0] addr_selector3_1173;
wire[15:0] addr_remain3_1173;
address_decode_4 decoder_3_1173 = address_decode_4(addr_selector2_73[5],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1173,addr_remain3_1173);


wire[15:0] addr_selector3_1174;
wire[15:0] addr_remain3_1174;
address_decode_4 decoder_3_1174 = address_decode_4(addr_selector2_73[6],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1174,addr_remain3_1174);


wire[15:0] addr_selector3_1175;
wire[15:0] addr_remain3_1175;
address_decode_4 decoder_3_1175 = address_decode_4(addr_selector2_73[7],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1175,addr_remain3_1175);


wire[15:0] addr_selector3_1176;
wire[15:0] addr_remain3_1176;
address_decode_4 decoder_3_1176 = address_decode_4(addr_selector2_73[8],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1176,addr_remain3_1176);


wire[15:0] addr_selector3_1177;
wire[15:0] addr_remain3_1177;
address_decode_4 decoder_3_1177 = address_decode_4(addr_selector2_73[9],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1177,addr_remain3_1177);


wire[15:0] addr_selector3_1178;
wire[15:0] addr_remain3_1178;
address_decode_4 decoder_3_1178 = address_decode_4(addr_selector2_73[10],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1178,addr_remain3_1178);


wire[15:0] addr_selector3_1179;
wire[15:0] addr_remain3_1179;
address_decode_4 decoder_3_1179 = address_decode_4(addr_selector2_73[11],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1179,addr_remain3_1179);


wire[15:0] addr_selector3_1180;
wire[15:0] addr_remain3_1180;
address_decode_4 decoder_3_1180 = address_decode_4(addr_selector2_73[12],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1180,addr_remain3_1180);


wire[15:0] addr_selector3_1181;
wire[15:0] addr_remain3_1181;
address_decode_4 decoder_3_1181 = address_decode_4(addr_selector2_73[13],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1181,addr_remain3_1181);


wire[15:0] addr_selector3_1182;
wire[15:0] addr_remain3_1182;
address_decode_4 decoder_3_1182 = address_decode_4(addr_selector2_73[14],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1182,addr_remain3_1182);


wire[15:0] addr_selector3_1183;
wire[15:0] addr_remain3_1183;
address_decode_4 decoder_3_1183 = address_decode_4(addr_selector2_73[15],addr_remain2_73[15:0],addr_remain2_73,addr_selector3_1183,addr_remain3_1183);


wire[15:0] addr_selector3_1184;
wire[15:0] addr_remain3_1184;
address_decode_4 decoder_3_1184 = address_decode_4(addr_selector2_74[0],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1184,addr_remain3_1184);


wire[15:0] addr_selector3_1185;
wire[15:0] addr_remain3_1185;
address_decode_4 decoder_3_1185 = address_decode_4(addr_selector2_74[1],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1185,addr_remain3_1185);


wire[15:0] addr_selector3_1186;
wire[15:0] addr_remain3_1186;
address_decode_4 decoder_3_1186 = address_decode_4(addr_selector2_74[2],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1186,addr_remain3_1186);


wire[15:0] addr_selector3_1187;
wire[15:0] addr_remain3_1187;
address_decode_4 decoder_3_1187 = address_decode_4(addr_selector2_74[3],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1187,addr_remain3_1187);


wire[15:0] addr_selector3_1188;
wire[15:0] addr_remain3_1188;
address_decode_4 decoder_3_1188 = address_decode_4(addr_selector2_74[4],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1188,addr_remain3_1188);


wire[15:0] addr_selector3_1189;
wire[15:0] addr_remain3_1189;
address_decode_4 decoder_3_1189 = address_decode_4(addr_selector2_74[5],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1189,addr_remain3_1189);


wire[15:0] addr_selector3_1190;
wire[15:0] addr_remain3_1190;
address_decode_4 decoder_3_1190 = address_decode_4(addr_selector2_74[6],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1190,addr_remain3_1190);


wire[15:0] addr_selector3_1191;
wire[15:0] addr_remain3_1191;
address_decode_4 decoder_3_1191 = address_decode_4(addr_selector2_74[7],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1191,addr_remain3_1191);


wire[15:0] addr_selector3_1192;
wire[15:0] addr_remain3_1192;
address_decode_4 decoder_3_1192 = address_decode_4(addr_selector2_74[8],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1192,addr_remain3_1192);


wire[15:0] addr_selector3_1193;
wire[15:0] addr_remain3_1193;
address_decode_4 decoder_3_1193 = address_decode_4(addr_selector2_74[9],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1193,addr_remain3_1193);


wire[15:0] addr_selector3_1194;
wire[15:0] addr_remain3_1194;
address_decode_4 decoder_3_1194 = address_decode_4(addr_selector2_74[10],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1194,addr_remain3_1194);


wire[15:0] addr_selector3_1195;
wire[15:0] addr_remain3_1195;
address_decode_4 decoder_3_1195 = address_decode_4(addr_selector2_74[11],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1195,addr_remain3_1195);


wire[15:0] addr_selector3_1196;
wire[15:0] addr_remain3_1196;
address_decode_4 decoder_3_1196 = address_decode_4(addr_selector2_74[12],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1196,addr_remain3_1196);


wire[15:0] addr_selector3_1197;
wire[15:0] addr_remain3_1197;
address_decode_4 decoder_3_1197 = address_decode_4(addr_selector2_74[13],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1197,addr_remain3_1197);


wire[15:0] addr_selector3_1198;
wire[15:0] addr_remain3_1198;
address_decode_4 decoder_3_1198 = address_decode_4(addr_selector2_74[14],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1198,addr_remain3_1198);


wire[15:0] addr_selector3_1199;
wire[15:0] addr_remain3_1199;
address_decode_4 decoder_3_1199 = address_decode_4(addr_selector2_74[15],addr_remain2_74[15:0],addr_remain2_74,addr_selector3_1199,addr_remain3_1199);


wire[15:0] addr_selector3_1200;
wire[15:0] addr_remain3_1200;
address_decode_4 decoder_3_1200 = address_decode_4(addr_selector2_75[0],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1200,addr_remain3_1200);


wire[15:0] addr_selector3_1201;
wire[15:0] addr_remain3_1201;
address_decode_4 decoder_3_1201 = address_decode_4(addr_selector2_75[1],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1201,addr_remain3_1201);


wire[15:0] addr_selector3_1202;
wire[15:0] addr_remain3_1202;
address_decode_4 decoder_3_1202 = address_decode_4(addr_selector2_75[2],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1202,addr_remain3_1202);


wire[15:0] addr_selector3_1203;
wire[15:0] addr_remain3_1203;
address_decode_4 decoder_3_1203 = address_decode_4(addr_selector2_75[3],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1203,addr_remain3_1203);


wire[15:0] addr_selector3_1204;
wire[15:0] addr_remain3_1204;
address_decode_4 decoder_3_1204 = address_decode_4(addr_selector2_75[4],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1204,addr_remain3_1204);


wire[15:0] addr_selector3_1205;
wire[15:0] addr_remain3_1205;
address_decode_4 decoder_3_1205 = address_decode_4(addr_selector2_75[5],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1205,addr_remain3_1205);


wire[15:0] addr_selector3_1206;
wire[15:0] addr_remain3_1206;
address_decode_4 decoder_3_1206 = address_decode_4(addr_selector2_75[6],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1206,addr_remain3_1206);


wire[15:0] addr_selector3_1207;
wire[15:0] addr_remain3_1207;
address_decode_4 decoder_3_1207 = address_decode_4(addr_selector2_75[7],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1207,addr_remain3_1207);


wire[15:0] addr_selector3_1208;
wire[15:0] addr_remain3_1208;
address_decode_4 decoder_3_1208 = address_decode_4(addr_selector2_75[8],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1208,addr_remain3_1208);


wire[15:0] addr_selector3_1209;
wire[15:0] addr_remain3_1209;
address_decode_4 decoder_3_1209 = address_decode_4(addr_selector2_75[9],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1209,addr_remain3_1209);


wire[15:0] addr_selector3_1210;
wire[15:0] addr_remain3_1210;
address_decode_4 decoder_3_1210 = address_decode_4(addr_selector2_75[10],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1210,addr_remain3_1210);


wire[15:0] addr_selector3_1211;
wire[15:0] addr_remain3_1211;
address_decode_4 decoder_3_1211 = address_decode_4(addr_selector2_75[11],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1211,addr_remain3_1211);


wire[15:0] addr_selector3_1212;
wire[15:0] addr_remain3_1212;
address_decode_4 decoder_3_1212 = address_decode_4(addr_selector2_75[12],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1212,addr_remain3_1212);


wire[15:0] addr_selector3_1213;
wire[15:0] addr_remain3_1213;
address_decode_4 decoder_3_1213 = address_decode_4(addr_selector2_75[13],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1213,addr_remain3_1213);


wire[15:0] addr_selector3_1214;
wire[15:0] addr_remain3_1214;
address_decode_4 decoder_3_1214 = address_decode_4(addr_selector2_75[14],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1214,addr_remain3_1214);


wire[15:0] addr_selector3_1215;
wire[15:0] addr_remain3_1215;
address_decode_4 decoder_3_1215 = address_decode_4(addr_selector2_75[15],addr_remain2_75[15:0],addr_remain2_75,addr_selector3_1215,addr_remain3_1215);


wire[15:0] addr_selector3_1216;
wire[15:0] addr_remain3_1216;
address_decode_4 decoder_3_1216 = address_decode_4(addr_selector2_76[0],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1216,addr_remain3_1216);


wire[15:0] addr_selector3_1217;
wire[15:0] addr_remain3_1217;
address_decode_4 decoder_3_1217 = address_decode_4(addr_selector2_76[1],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1217,addr_remain3_1217);


wire[15:0] addr_selector3_1218;
wire[15:0] addr_remain3_1218;
address_decode_4 decoder_3_1218 = address_decode_4(addr_selector2_76[2],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1218,addr_remain3_1218);


wire[15:0] addr_selector3_1219;
wire[15:0] addr_remain3_1219;
address_decode_4 decoder_3_1219 = address_decode_4(addr_selector2_76[3],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1219,addr_remain3_1219);


wire[15:0] addr_selector3_1220;
wire[15:0] addr_remain3_1220;
address_decode_4 decoder_3_1220 = address_decode_4(addr_selector2_76[4],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1220,addr_remain3_1220);


wire[15:0] addr_selector3_1221;
wire[15:0] addr_remain3_1221;
address_decode_4 decoder_3_1221 = address_decode_4(addr_selector2_76[5],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1221,addr_remain3_1221);


wire[15:0] addr_selector3_1222;
wire[15:0] addr_remain3_1222;
address_decode_4 decoder_3_1222 = address_decode_4(addr_selector2_76[6],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1222,addr_remain3_1222);


wire[15:0] addr_selector3_1223;
wire[15:0] addr_remain3_1223;
address_decode_4 decoder_3_1223 = address_decode_4(addr_selector2_76[7],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1223,addr_remain3_1223);


wire[15:0] addr_selector3_1224;
wire[15:0] addr_remain3_1224;
address_decode_4 decoder_3_1224 = address_decode_4(addr_selector2_76[8],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1224,addr_remain3_1224);


wire[15:0] addr_selector3_1225;
wire[15:0] addr_remain3_1225;
address_decode_4 decoder_3_1225 = address_decode_4(addr_selector2_76[9],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1225,addr_remain3_1225);


wire[15:0] addr_selector3_1226;
wire[15:0] addr_remain3_1226;
address_decode_4 decoder_3_1226 = address_decode_4(addr_selector2_76[10],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1226,addr_remain3_1226);


wire[15:0] addr_selector3_1227;
wire[15:0] addr_remain3_1227;
address_decode_4 decoder_3_1227 = address_decode_4(addr_selector2_76[11],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1227,addr_remain3_1227);


wire[15:0] addr_selector3_1228;
wire[15:0] addr_remain3_1228;
address_decode_4 decoder_3_1228 = address_decode_4(addr_selector2_76[12],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1228,addr_remain3_1228);


wire[15:0] addr_selector3_1229;
wire[15:0] addr_remain3_1229;
address_decode_4 decoder_3_1229 = address_decode_4(addr_selector2_76[13],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1229,addr_remain3_1229);


wire[15:0] addr_selector3_1230;
wire[15:0] addr_remain3_1230;
address_decode_4 decoder_3_1230 = address_decode_4(addr_selector2_76[14],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1230,addr_remain3_1230);


wire[15:0] addr_selector3_1231;
wire[15:0] addr_remain3_1231;
address_decode_4 decoder_3_1231 = address_decode_4(addr_selector2_76[15],addr_remain2_76[15:0],addr_remain2_76,addr_selector3_1231,addr_remain3_1231);


wire[15:0] addr_selector3_1232;
wire[15:0] addr_remain3_1232;
address_decode_4 decoder_3_1232 = address_decode_4(addr_selector2_77[0],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1232,addr_remain3_1232);


wire[15:0] addr_selector3_1233;
wire[15:0] addr_remain3_1233;
address_decode_4 decoder_3_1233 = address_decode_4(addr_selector2_77[1],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1233,addr_remain3_1233);


wire[15:0] addr_selector3_1234;
wire[15:0] addr_remain3_1234;
address_decode_4 decoder_3_1234 = address_decode_4(addr_selector2_77[2],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1234,addr_remain3_1234);


wire[15:0] addr_selector3_1235;
wire[15:0] addr_remain3_1235;
address_decode_4 decoder_3_1235 = address_decode_4(addr_selector2_77[3],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1235,addr_remain3_1235);


wire[15:0] addr_selector3_1236;
wire[15:0] addr_remain3_1236;
address_decode_4 decoder_3_1236 = address_decode_4(addr_selector2_77[4],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1236,addr_remain3_1236);


wire[15:0] addr_selector3_1237;
wire[15:0] addr_remain3_1237;
address_decode_4 decoder_3_1237 = address_decode_4(addr_selector2_77[5],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1237,addr_remain3_1237);


wire[15:0] addr_selector3_1238;
wire[15:0] addr_remain3_1238;
address_decode_4 decoder_3_1238 = address_decode_4(addr_selector2_77[6],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1238,addr_remain3_1238);


wire[15:0] addr_selector3_1239;
wire[15:0] addr_remain3_1239;
address_decode_4 decoder_3_1239 = address_decode_4(addr_selector2_77[7],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1239,addr_remain3_1239);


wire[15:0] addr_selector3_1240;
wire[15:0] addr_remain3_1240;
address_decode_4 decoder_3_1240 = address_decode_4(addr_selector2_77[8],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1240,addr_remain3_1240);


wire[15:0] addr_selector3_1241;
wire[15:0] addr_remain3_1241;
address_decode_4 decoder_3_1241 = address_decode_4(addr_selector2_77[9],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1241,addr_remain3_1241);


wire[15:0] addr_selector3_1242;
wire[15:0] addr_remain3_1242;
address_decode_4 decoder_3_1242 = address_decode_4(addr_selector2_77[10],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1242,addr_remain3_1242);


wire[15:0] addr_selector3_1243;
wire[15:0] addr_remain3_1243;
address_decode_4 decoder_3_1243 = address_decode_4(addr_selector2_77[11],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1243,addr_remain3_1243);


wire[15:0] addr_selector3_1244;
wire[15:0] addr_remain3_1244;
address_decode_4 decoder_3_1244 = address_decode_4(addr_selector2_77[12],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1244,addr_remain3_1244);


wire[15:0] addr_selector3_1245;
wire[15:0] addr_remain3_1245;
address_decode_4 decoder_3_1245 = address_decode_4(addr_selector2_77[13],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1245,addr_remain3_1245);


wire[15:0] addr_selector3_1246;
wire[15:0] addr_remain3_1246;
address_decode_4 decoder_3_1246 = address_decode_4(addr_selector2_77[14],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1246,addr_remain3_1246);


wire[15:0] addr_selector3_1247;
wire[15:0] addr_remain3_1247;
address_decode_4 decoder_3_1247 = address_decode_4(addr_selector2_77[15],addr_remain2_77[15:0],addr_remain2_77,addr_selector3_1247,addr_remain3_1247);


wire[15:0] addr_selector3_1248;
wire[15:0] addr_remain3_1248;
address_decode_4 decoder_3_1248 = address_decode_4(addr_selector2_78[0],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1248,addr_remain3_1248);


wire[15:0] addr_selector3_1249;
wire[15:0] addr_remain3_1249;
address_decode_4 decoder_3_1249 = address_decode_4(addr_selector2_78[1],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1249,addr_remain3_1249);


wire[15:0] addr_selector3_1250;
wire[15:0] addr_remain3_1250;
address_decode_4 decoder_3_1250 = address_decode_4(addr_selector2_78[2],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1250,addr_remain3_1250);


wire[15:0] addr_selector3_1251;
wire[15:0] addr_remain3_1251;
address_decode_4 decoder_3_1251 = address_decode_4(addr_selector2_78[3],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1251,addr_remain3_1251);


wire[15:0] addr_selector3_1252;
wire[15:0] addr_remain3_1252;
address_decode_4 decoder_3_1252 = address_decode_4(addr_selector2_78[4],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1252,addr_remain3_1252);


wire[15:0] addr_selector3_1253;
wire[15:0] addr_remain3_1253;
address_decode_4 decoder_3_1253 = address_decode_4(addr_selector2_78[5],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1253,addr_remain3_1253);


wire[15:0] addr_selector3_1254;
wire[15:0] addr_remain3_1254;
address_decode_4 decoder_3_1254 = address_decode_4(addr_selector2_78[6],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1254,addr_remain3_1254);


wire[15:0] addr_selector3_1255;
wire[15:0] addr_remain3_1255;
address_decode_4 decoder_3_1255 = address_decode_4(addr_selector2_78[7],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1255,addr_remain3_1255);


wire[15:0] addr_selector3_1256;
wire[15:0] addr_remain3_1256;
address_decode_4 decoder_3_1256 = address_decode_4(addr_selector2_78[8],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1256,addr_remain3_1256);


wire[15:0] addr_selector3_1257;
wire[15:0] addr_remain3_1257;
address_decode_4 decoder_3_1257 = address_decode_4(addr_selector2_78[9],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1257,addr_remain3_1257);


wire[15:0] addr_selector3_1258;
wire[15:0] addr_remain3_1258;
address_decode_4 decoder_3_1258 = address_decode_4(addr_selector2_78[10],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1258,addr_remain3_1258);


wire[15:0] addr_selector3_1259;
wire[15:0] addr_remain3_1259;
address_decode_4 decoder_3_1259 = address_decode_4(addr_selector2_78[11],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1259,addr_remain3_1259);


wire[15:0] addr_selector3_1260;
wire[15:0] addr_remain3_1260;
address_decode_4 decoder_3_1260 = address_decode_4(addr_selector2_78[12],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1260,addr_remain3_1260);


wire[15:0] addr_selector3_1261;
wire[15:0] addr_remain3_1261;
address_decode_4 decoder_3_1261 = address_decode_4(addr_selector2_78[13],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1261,addr_remain3_1261);


wire[15:0] addr_selector3_1262;
wire[15:0] addr_remain3_1262;
address_decode_4 decoder_3_1262 = address_decode_4(addr_selector2_78[14],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1262,addr_remain3_1262);


wire[15:0] addr_selector3_1263;
wire[15:0] addr_remain3_1263;
address_decode_4 decoder_3_1263 = address_decode_4(addr_selector2_78[15],addr_remain2_78[15:0],addr_remain2_78,addr_selector3_1263,addr_remain3_1263);


wire[15:0] addr_selector3_1264;
wire[15:0] addr_remain3_1264;
address_decode_4 decoder_3_1264 = address_decode_4(addr_selector2_79[0],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1264,addr_remain3_1264);


wire[15:0] addr_selector3_1265;
wire[15:0] addr_remain3_1265;
address_decode_4 decoder_3_1265 = address_decode_4(addr_selector2_79[1],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1265,addr_remain3_1265);


wire[15:0] addr_selector3_1266;
wire[15:0] addr_remain3_1266;
address_decode_4 decoder_3_1266 = address_decode_4(addr_selector2_79[2],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1266,addr_remain3_1266);


wire[15:0] addr_selector3_1267;
wire[15:0] addr_remain3_1267;
address_decode_4 decoder_3_1267 = address_decode_4(addr_selector2_79[3],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1267,addr_remain3_1267);


wire[15:0] addr_selector3_1268;
wire[15:0] addr_remain3_1268;
address_decode_4 decoder_3_1268 = address_decode_4(addr_selector2_79[4],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1268,addr_remain3_1268);


wire[15:0] addr_selector3_1269;
wire[15:0] addr_remain3_1269;
address_decode_4 decoder_3_1269 = address_decode_4(addr_selector2_79[5],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1269,addr_remain3_1269);


wire[15:0] addr_selector3_1270;
wire[15:0] addr_remain3_1270;
address_decode_4 decoder_3_1270 = address_decode_4(addr_selector2_79[6],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1270,addr_remain3_1270);


wire[15:0] addr_selector3_1271;
wire[15:0] addr_remain3_1271;
address_decode_4 decoder_3_1271 = address_decode_4(addr_selector2_79[7],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1271,addr_remain3_1271);


wire[15:0] addr_selector3_1272;
wire[15:0] addr_remain3_1272;
address_decode_4 decoder_3_1272 = address_decode_4(addr_selector2_79[8],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1272,addr_remain3_1272);


wire[15:0] addr_selector3_1273;
wire[15:0] addr_remain3_1273;
address_decode_4 decoder_3_1273 = address_decode_4(addr_selector2_79[9],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1273,addr_remain3_1273);


wire[15:0] addr_selector3_1274;
wire[15:0] addr_remain3_1274;
address_decode_4 decoder_3_1274 = address_decode_4(addr_selector2_79[10],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1274,addr_remain3_1274);


wire[15:0] addr_selector3_1275;
wire[15:0] addr_remain3_1275;
address_decode_4 decoder_3_1275 = address_decode_4(addr_selector2_79[11],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1275,addr_remain3_1275);


wire[15:0] addr_selector3_1276;
wire[15:0] addr_remain3_1276;
address_decode_4 decoder_3_1276 = address_decode_4(addr_selector2_79[12],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1276,addr_remain3_1276);


wire[15:0] addr_selector3_1277;
wire[15:0] addr_remain3_1277;
address_decode_4 decoder_3_1277 = address_decode_4(addr_selector2_79[13],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1277,addr_remain3_1277);


wire[15:0] addr_selector3_1278;
wire[15:0] addr_remain3_1278;
address_decode_4 decoder_3_1278 = address_decode_4(addr_selector2_79[14],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1278,addr_remain3_1278);


wire[15:0] addr_selector3_1279;
wire[15:0] addr_remain3_1279;
address_decode_4 decoder_3_1279 = address_decode_4(addr_selector2_79[15],addr_remain2_79[15:0],addr_remain2_79,addr_selector3_1279,addr_remain3_1279);


wire[15:0] addr_selector3_1280;
wire[15:0] addr_remain3_1280;
address_decode_4 decoder_3_1280 = address_decode_4(addr_selector2_80[0],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1280,addr_remain3_1280);


wire[15:0] addr_selector3_1281;
wire[15:0] addr_remain3_1281;
address_decode_4 decoder_3_1281 = address_decode_4(addr_selector2_80[1],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1281,addr_remain3_1281);


wire[15:0] addr_selector3_1282;
wire[15:0] addr_remain3_1282;
address_decode_4 decoder_3_1282 = address_decode_4(addr_selector2_80[2],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1282,addr_remain3_1282);


wire[15:0] addr_selector3_1283;
wire[15:0] addr_remain3_1283;
address_decode_4 decoder_3_1283 = address_decode_4(addr_selector2_80[3],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1283,addr_remain3_1283);


wire[15:0] addr_selector3_1284;
wire[15:0] addr_remain3_1284;
address_decode_4 decoder_3_1284 = address_decode_4(addr_selector2_80[4],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1284,addr_remain3_1284);


wire[15:0] addr_selector3_1285;
wire[15:0] addr_remain3_1285;
address_decode_4 decoder_3_1285 = address_decode_4(addr_selector2_80[5],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1285,addr_remain3_1285);


wire[15:0] addr_selector3_1286;
wire[15:0] addr_remain3_1286;
address_decode_4 decoder_3_1286 = address_decode_4(addr_selector2_80[6],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1286,addr_remain3_1286);


wire[15:0] addr_selector3_1287;
wire[15:0] addr_remain3_1287;
address_decode_4 decoder_3_1287 = address_decode_4(addr_selector2_80[7],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1287,addr_remain3_1287);


wire[15:0] addr_selector3_1288;
wire[15:0] addr_remain3_1288;
address_decode_4 decoder_3_1288 = address_decode_4(addr_selector2_80[8],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1288,addr_remain3_1288);


wire[15:0] addr_selector3_1289;
wire[15:0] addr_remain3_1289;
address_decode_4 decoder_3_1289 = address_decode_4(addr_selector2_80[9],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1289,addr_remain3_1289);


wire[15:0] addr_selector3_1290;
wire[15:0] addr_remain3_1290;
address_decode_4 decoder_3_1290 = address_decode_4(addr_selector2_80[10],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1290,addr_remain3_1290);


wire[15:0] addr_selector3_1291;
wire[15:0] addr_remain3_1291;
address_decode_4 decoder_3_1291 = address_decode_4(addr_selector2_80[11],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1291,addr_remain3_1291);


wire[15:0] addr_selector3_1292;
wire[15:0] addr_remain3_1292;
address_decode_4 decoder_3_1292 = address_decode_4(addr_selector2_80[12],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1292,addr_remain3_1292);


wire[15:0] addr_selector3_1293;
wire[15:0] addr_remain3_1293;
address_decode_4 decoder_3_1293 = address_decode_4(addr_selector2_80[13],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1293,addr_remain3_1293);


wire[15:0] addr_selector3_1294;
wire[15:0] addr_remain3_1294;
address_decode_4 decoder_3_1294 = address_decode_4(addr_selector2_80[14],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1294,addr_remain3_1294);


wire[15:0] addr_selector3_1295;
wire[15:0] addr_remain3_1295;
address_decode_4 decoder_3_1295 = address_decode_4(addr_selector2_80[15],addr_remain2_80[15:0],addr_remain2_80,addr_selector3_1295,addr_remain3_1295);


wire[15:0] addr_selector3_1296;
wire[15:0] addr_remain3_1296;
address_decode_4 decoder_3_1296 = address_decode_4(addr_selector2_81[0],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1296,addr_remain3_1296);


wire[15:0] addr_selector3_1297;
wire[15:0] addr_remain3_1297;
address_decode_4 decoder_3_1297 = address_decode_4(addr_selector2_81[1],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1297,addr_remain3_1297);


wire[15:0] addr_selector3_1298;
wire[15:0] addr_remain3_1298;
address_decode_4 decoder_3_1298 = address_decode_4(addr_selector2_81[2],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1298,addr_remain3_1298);


wire[15:0] addr_selector3_1299;
wire[15:0] addr_remain3_1299;
address_decode_4 decoder_3_1299 = address_decode_4(addr_selector2_81[3],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1299,addr_remain3_1299);


wire[15:0] addr_selector3_1300;
wire[15:0] addr_remain3_1300;
address_decode_4 decoder_3_1300 = address_decode_4(addr_selector2_81[4],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1300,addr_remain3_1300);


wire[15:0] addr_selector3_1301;
wire[15:0] addr_remain3_1301;
address_decode_4 decoder_3_1301 = address_decode_4(addr_selector2_81[5],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1301,addr_remain3_1301);


wire[15:0] addr_selector3_1302;
wire[15:0] addr_remain3_1302;
address_decode_4 decoder_3_1302 = address_decode_4(addr_selector2_81[6],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1302,addr_remain3_1302);


wire[15:0] addr_selector3_1303;
wire[15:0] addr_remain3_1303;
address_decode_4 decoder_3_1303 = address_decode_4(addr_selector2_81[7],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1303,addr_remain3_1303);


wire[15:0] addr_selector3_1304;
wire[15:0] addr_remain3_1304;
address_decode_4 decoder_3_1304 = address_decode_4(addr_selector2_81[8],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1304,addr_remain3_1304);


wire[15:0] addr_selector3_1305;
wire[15:0] addr_remain3_1305;
address_decode_4 decoder_3_1305 = address_decode_4(addr_selector2_81[9],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1305,addr_remain3_1305);


wire[15:0] addr_selector3_1306;
wire[15:0] addr_remain3_1306;
address_decode_4 decoder_3_1306 = address_decode_4(addr_selector2_81[10],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1306,addr_remain3_1306);


wire[15:0] addr_selector3_1307;
wire[15:0] addr_remain3_1307;
address_decode_4 decoder_3_1307 = address_decode_4(addr_selector2_81[11],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1307,addr_remain3_1307);


wire[15:0] addr_selector3_1308;
wire[15:0] addr_remain3_1308;
address_decode_4 decoder_3_1308 = address_decode_4(addr_selector2_81[12],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1308,addr_remain3_1308);


wire[15:0] addr_selector3_1309;
wire[15:0] addr_remain3_1309;
address_decode_4 decoder_3_1309 = address_decode_4(addr_selector2_81[13],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1309,addr_remain3_1309);


wire[15:0] addr_selector3_1310;
wire[15:0] addr_remain3_1310;
address_decode_4 decoder_3_1310 = address_decode_4(addr_selector2_81[14],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1310,addr_remain3_1310);


wire[15:0] addr_selector3_1311;
wire[15:0] addr_remain3_1311;
address_decode_4 decoder_3_1311 = address_decode_4(addr_selector2_81[15],addr_remain2_81[15:0],addr_remain2_81,addr_selector3_1311,addr_remain3_1311);


wire[15:0] addr_selector3_1312;
wire[15:0] addr_remain3_1312;
address_decode_4 decoder_3_1312 = address_decode_4(addr_selector2_82[0],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1312,addr_remain3_1312);


wire[15:0] addr_selector3_1313;
wire[15:0] addr_remain3_1313;
address_decode_4 decoder_3_1313 = address_decode_4(addr_selector2_82[1],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1313,addr_remain3_1313);


wire[15:0] addr_selector3_1314;
wire[15:0] addr_remain3_1314;
address_decode_4 decoder_3_1314 = address_decode_4(addr_selector2_82[2],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1314,addr_remain3_1314);


wire[15:0] addr_selector3_1315;
wire[15:0] addr_remain3_1315;
address_decode_4 decoder_3_1315 = address_decode_4(addr_selector2_82[3],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1315,addr_remain3_1315);


wire[15:0] addr_selector3_1316;
wire[15:0] addr_remain3_1316;
address_decode_4 decoder_3_1316 = address_decode_4(addr_selector2_82[4],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1316,addr_remain3_1316);


wire[15:0] addr_selector3_1317;
wire[15:0] addr_remain3_1317;
address_decode_4 decoder_3_1317 = address_decode_4(addr_selector2_82[5],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1317,addr_remain3_1317);


wire[15:0] addr_selector3_1318;
wire[15:0] addr_remain3_1318;
address_decode_4 decoder_3_1318 = address_decode_4(addr_selector2_82[6],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1318,addr_remain3_1318);


wire[15:0] addr_selector3_1319;
wire[15:0] addr_remain3_1319;
address_decode_4 decoder_3_1319 = address_decode_4(addr_selector2_82[7],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1319,addr_remain3_1319);


wire[15:0] addr_selector3_1320;
wire[15:0] addr_remain3_1320;
address_decode_4 decoder_3_1320 = address_decode_4(addr_selector2_82[8],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1320,addr_remain3_1320);


wire[15:0] addr_selector3_1321;
wire[15:0] addr_remain3_1321;
address_decode_4 decoder_3_1321 = address_decode_4(addr_selector2_82[9],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1321,addr_remain3_1321);


wire[15:0] addr_selector3_1322;
wire[15:0] addr_remain3_1322;
address_decode_4 decoder_3_1322 = address_decode_4(addr_selector2_82[10],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1322,addr_remain3_1322);


wire[15:0] addr_selector3_1323;
wire[15:0] addr_remain3_1323;
address_decode_4 decoder_3_1323 = address_decode_4(addr_selector2_82[11],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1323,addr_remain3_1323);


wire[15:0] addr_selector3_1324;
wire[15:0] addr_remain3_1324;
address_decode_4 decoder_3_1324 = address_decode_4(addr_selector2_82[12],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1324,addr_remain3_1324);


wire[15:0] addr_selector3_1325;
wire[15:0] addr_remain3_1325;
address_decode_4 decoder_3_1325 = address_decode_4(addr_selector2_82[13],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1325,addr_remain3_1325);


wire[15:0] addr_selector3_1326;
wire[15:0] addr_remain3_1326;
address_decode_4 decoder_3_1326 = address_decode_4(addr_selector2_82[14],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1326,addr_remain3_1326);


wire[15:0] addr_selector3_1327;
wire[15:0] addr_remain3_1327;
address_decode_4 decoder_3_1327 = address_decode_4(addr_selector2_82[15],addr_remain2_82[15:0],addr_remain2_82,addr_selector3_1327,addr_remain3_1327);


wire[15:0] addr_selector3_1328;
wire[15:0] addr_remain3_1328;
address_decode_4 decoder_3_1328 = address_decode_4(addr_selector2_83[0],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1328,addr_remain3_1328);


wire[15:0] addr_selector3_1329;
wire[15:0] addr_remain3_1329;
address_decode_4 decoder_3_1329 = address_decode_4(addr_selector2_83[1],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1329,addr_remain3_1329);


wire[15:0] addr_selector3_1330;
wire[15:0] addr_remain3_1330;
address_decode_4 decoder_3_1330 = address_decode_4(addr_selector2_83[2],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1330,addr_remain3_1330);


wire[15:0] addr_selector3_1331;
wire[15:0] addr_remain3_1331;
address_decode_4 decoder_3_1331 = address_decode_4(addr_selector2_83[3],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1331,addr_remain3_1331);


wire[15:0] addr_selector3_1332;
wire[15:0] addr_remain3_1332;
address_decode_4 decoder_3_1332 = address_decode_4(addr_selector2_83[4],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1332,addr_remain3_1332);


wire[15:0] addr_selector3_1333;
wire[15:0] addr_remain3_1333;
address_decode_4 decoder_3_1333 = address_decode_4(addr_selector2_83[5],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1333,addr_remain3_1333);


wire[15:0] addr_selector3_1334;
wire[15:0] addr_remain3_1334;
address_decode_4 decoder_3_1334 = address_decode_4(addr_selector2_83[6],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1334,addr_remain3_1334);


wire[15:0] addr_selector3_1335;
wire[15:0] addr_remain3_1335;
address_decode_4 decoder_3_1335 = address_decode_4(addr_selector2_83[7],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1335,addr_remain3_1335);


wire[15:0] addr_selector3_1336;
wire[15:0] addr_remain3_1336;
address_decode_4 decoder_3_1336 = address_decode_4(addr_selector2_83[8],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1336,addr_remain3_1336);


wire[15:0] addr_selector3_1337;
wire[15:0] addr_remain3_1337;
address_decode_4 decoder_3_1337 = address_decode_4(addr_selector2_83[9],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1337,addr_remain3_1337);


wire[15:0] addr_selector3_1338;
wire[15:0] addr_remain3_1338;
address_decode_4 decoder_3_1338 = address_decode_4(addr_selector2_83[10],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1338,addr_remain3_1338);


wire[15:0] addr_selector3_1339;
wire[15:0] addr_remain3_1339;
address_decode_4 decoder_3_1339 = address_decode_4(addr_selector2_83[11],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1339,addr_remain3_1339);


wire[15:0] addr_selector3_1340;
wire[15:0] addr_remain3_1340;
address_decode_4 decoder_3_1340 = address_decode_4(addr_selector2_83[12],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1340,addr_remain3_1340);


wire[15:0] addr_selector3_1341;
wire[15:0] addr_remain3_1341;
address_decode_4 decoder_3_1341 = address_decode_4(addr_selector2_83[13],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1341,addr_remain3_1341);


wire[15:0] addr_selector3_1342;
wire[15:0] addr_remain3_1342;
address_decode_4 decoder_3_1342 = address_decode_4(addr_selector2_83[14],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1342,addr_remain3_1342);


wire[15:0] addr_selector3_1343;
wire[15:0] addr_remain3_1343;
address_decode_4 decoder_3_1343 = address_decode_4(addr_selector2_83[15],addr_remain2_83[15:0],addr_remain2_83,addr_selector3_1343,addr_remain3_1343);


wire[15:0] addr_selector3_1344;
wire[15:0] addr_remain3_1344;
address_decode_4 decoder_3_1344 = address_decode_4(addr_selector2_84[0],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1344,addr_remain3_1344);


wire[15:0] addr_selector3_1345;
wire[15:0] addr_remain3_1345;
address_decode_4 decoder_3_1345 = address_decode_4(addr_selector2_84[1],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1345,addr_remain3_1345);


wire[15:0] addr_selector3_1346;
wire[15:0] addr_remain3_1346;
address_decode_4 decoder_3_1346 = address_decode_4(addr_selector2_84[2],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1346,addr_remain3_1346);


wire[15:0] addr_selector3_1347;
wire[15:0] addr_remain3_1347;
address_decode_4 decoder_3_1347 = address_decode_4(addr_selector2_84[3],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1347,addr_remain3_1347);


wire[15:0] addr_selector3_1348;
wire[15:0] addr_remain3_1348;
address_decode_4 decoder_3_1348 = address_decode_4(addr_selector2_84[4],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1348,addr_remain3_1348);


wire[15:0] addr_selector3_1349;
wire[15:0] addr_remain3_1349;
address_decode_4 decoder_3_1349 = address_decode_4(addr_selector2_84[5],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1349,addr_remain3_1349);


wire[15:0] addr_selector3_1350;
wire[15:0] addr_remain3_1350;
address_decode_4 decoder_3_1350 = address_decode_4(addr_selector2_84[6],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1350,addr_remain3_1350);


wire[15:0] addr_selector3_1351;
wire[15:0] addr_remain3_1351;
address_decode_4 decoder_3_1351 = address_decode_4(addr_selector2_84[7],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1351,addr_remain3_1351);


wire[15:0] addr_selector3_1352;
wire[15:0] addr_remain3_1352;
address_decode_4 decoder_3_1352 = address_decode_4(addr_selector2_84[8],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1352,addr_remain3_1352);


wire[15:0] addr_selector3_1353;
wire[15:0] addr_remain3_1353;
address_decode_4 decoder_3_1353 = address_decode_4(addr_selector2_84[9],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1353,addr_remain3_1353);


wire[15:0] addr_selector3_1354;
wire[15:0] addr_remain3_1354;
address_decode_4 decoder_3_1354 = address_decode_4(addr_selector2_84[10],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1354,addr_remain3_1354);


wire[15:0] addr_selector3_1355;
wire[15:0] addr_remain3_1355;
address_decode_4 decoder_3_1355 = address_decode_4(addr_selector2_84[11],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1355,addr_remain3_1355);


wire[15:0] addr_selector3_1356;
wire[15:0] addr_remain3_1356;
address_decode_4 decoder_3_1356 = address_decode_4(addr_selector2_84[12],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1356,addr_remain3_1356);


wire[15:0] addr_selector3_1357;
wire[15:0] addr_remain3_1357;
address_decode_4 decoder_3_1357 = address_decode_4(addr_selector2_84[13],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1357,addr_remain3_1357);


wire[15:0] addr_selector3_1358;
wire[15:0] addr_remain3_1358;
address_decode_4 decoder_3_1358 = address_decode_4(addr_selector2_84[14],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1358,addr_remain3_1358);


wire[15:0] addr_selector3_1359;
wire[15:0] addr_remain3_1359;
address_decode_4 decoder_3_1359 = address_decode_4(addr_selector2_84[15],addr_remain2_84[15:0],addr_remain2_84,addr_selector3_1359,addr_remain3_1359);


wire[15:0] addr_selector3_1360;
wire[15:0] addr_remain3_1360;
address_decode_4 decoder_3_1360 = address_decode_4(addr_selector2_85[0],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1360,addr_remain3_1360);


wire[15:0] addr_selector3_1361;
wire[15:0] addr_remain3_1361;
address_decode_4 decoder_3_1361 = address_decode_4(addr_selector2_85[1],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1361,addr_remain3_1361);


wire[15:0] addr_selector3_1362;
wire[15:0] addr_remain3_1362;
address_decode_4 decoder_3_1362 = address_decode_4(addr_selector2_85[2],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1362,addr_remain3_1362);


wire[15:0] addr_selector3_1363;
wire[15:0] addr_remain3_1363;
address_decode_4 decoder_3_1363 = address_decode_4(addr_selector2_85[3],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1363,addr_remain3_1363);


wire[15:0] addr_selector3_1364;
wire[15:0] addr_remain3_1364;
address_decode_4 decoder_3_1364 = address_decode_4(addr_selector2_85[4],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1364,addr_remain3_1364);


wire[15:0] addr_selector3_1365;
wire[15:0] addr_remain3_1365;
address_decode_4 decoder_3_1365 = address_decode_4(addr_selector2_85[5],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1365,addr_remain3_1365);


wire[15:0] addr_selector3_1366;
wire[15:0] addr_remain3_1366;
address_decode_4 decoder_3_1366 = address_decode_4(addr_selector2_85[6],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1366,addr_remain3_1366);


wire[15:0] addr_selector3_1367;
wire[15:0] addr_remain3_1367;
address_decode_4 decoder_3_1367 = address_decode_4(addr_selector2_85[7],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1367,addr_remain3_1367);


wire[15:0] addr_selector3_1368;
wire[15:0] addr_remain3_1368;
address_decode_4 decoder_3_1368 = address_decode_4(addr_selector2_85[8],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1368,addr_remain3_1368);


wire[15:0] addr_selector3_1369;
wire[15:0] addr_remain3_1369;
address_decode_4 decoder_3_1369 = address_decode_4(addr_selector2_85[9],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1369,addr_remain3_1369);


wire[15:0] addr_selector3_1370;
wire[15:0] addr_remain3_1370;
address_decode_4 decoder_3_1370 = address_decode_4(addr_selector2_85[10],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1370,addr_remain3_1370);


wire[15:0] addr_selector3_1371;
wire[15:0] addr_remain3_1371;
address_decode_4 decoder_3_1371 = address_decode_4(addr_selector2_85[11],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1371,addr_remain3_1371);


wire[15:0] addr_selector3_1372;
wire[15:0] addr_remain3_1372;
address_decode_4 decoder_3_1372 = address_decode_4(addr_selector2_85[12],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1372,addr_remain3_1372);


wire[15:0] addr_selector3_1373;
wire[15:0] addr_remain3_1373;
address_decode_4 decoder_3_1373 = address_decode_4(addr_selector2_85[13],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1373,addr_remain3_1373);


wire[15:0] addr_selector3_1374;
wire[15:0] addr_remain3_1374;
address_decode_4 decoder_3_1374 = address_decode_4(addr_selector2_85[14],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1374,addr_remain3_1374);


wire[15:0] addr_selector3_1375;
wire[15:0] addr_remain3_1375;
address_decode_4 decoder_3_1375 = address_decode_4(addr_selector2_85[15],addr_remain2_85[15:0],addr_remain2_85,addr_selector3_1375,addr_remain3_1375);


wire[15:0] addr_selector3_1376;
wire[15:0] addr_remain3_1376;
address_decode_4 decoder_3_1376 = address_decode_4(addr_selector2_86[0],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1376,addr_remain3_1376);


wire[15:0] addr_selector3_1377;
wire[15:0] addr_remain3_1377;
address_decode_4 decoder_3_1377 = address_decode_4(addr_selector2_86[1],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1377,addr_remain3_1377);


wire[15:0] addr_selector3_1378;
wire[15:0] addr_remain3_1378;
address_decode_4 decoder_3_1378 = address_decode_4(addr_selector2_86[2],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1378,addr_remain3_1378);


wire[15:0] addr_selector3_1379;
wire[15:0] addr_remain3_1379;
address_decode_4 decoder_3_1379 = address_decode_4(addr_selector2_86[3],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1379,addr_remain3_1379);


wire[15:0] addr_selector3_1380;
wire[15:0] addr_remain3_1380;
address_decode_4 decoder_3_1380 = address_decode_4(addr_selector2_86[4],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1380,addr_remain3_1380);


wire[15:0] addr_selector3_1381;
wire[15:0] addr_remain3_1381;
address_decode_4 decoder_3_1381 = address_decode_4(addr_selector2_86[5],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1381,addr_remain3_1381);


wire[15:0] addr_selector3_1382;
wire[15:0] addr_remain3_1382;
address_decode_4 decoder_3_1382 = address_decode_4(addr_selector2_86[6],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1382,addr_remain3_1382);


wire[15:0] addr_selector3_1383;
wire[15:0] addr_remain3_1383;
address_decode_4 decoder_3_1383 = address_decode_4(addr_selector2_86[7],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1383,addr_remain3_1383);


wire[15:0] addr_selector3_1384;
wire[15:0] addr_remain3_1384;
address_decode_4 decoder_3_1384 = address_decode_4(addr_selector2_86[8],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1384,addr_remain3_1384);


wire[15:0] addr_selector3_1385;
wire[15:0] addr_remain3_1385;
address_decode_4 decoder_3_1385 = address_decode_4(addr_selector2_86[9],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1385,addr_remain3_1385);


wire[15:0] addr_selector3_1386;
wire[15:0] addr_remain3_1386;
address_decode_4 decoder_3_1386 = address_decode_4(addr_selector2_86[10],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1386,addr_remain3_1386);


wire[15:0] addr_selector3_1387;
wire[15:0] addr_remain3_1387;
address_decode_4 decoder_3_1387 = address_decode_4(addr_selector2_86[11],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1387,addr_remain3_1387);


wire[15:0] addr_selector3_1388;
wire[15:0] addr_remain3_1388;
address_decode_4 decoder_3_1388 = address_decode_4(addr_selector2_86[12],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1388,addr_remain3_1388);


wire[15:0] addr_selector3_1389;
wire[15:0] addr_remain3_1389;
address_decode_4 decoder_3_1389 = address_decode_4(addr_selector2_86[13],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1389,addr_remain3_1389);


wire[15:0] addr_selector3_1390;
wire[15:0] addr_remain3_1390;
address_decode_4 decoder_3_1390 = address_decode_4(addr_selector2_86[14],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1390,addr_remain3_1390);


wire[15:0] addr_selector3_1391;
wire[15:0] addr_remain3_1391;
address_decode_4 decoder_3_1391 = address_decode_4(addr_selector2_86[15],addr_remain2_86[15:0],addr_remain2_86,addr_selector3_1391,addr_remain3_1391);


wire[15:0] addr_selector3_1392;
wire[15:0] addr_remain3_1392;
address_decode_4 decoder_3_1392 = address_decode_4(addr_selector2_87[0],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1392,addr_remain3_1392);


wire[15:0] addr_selector3_1393;
wire[15:0] addr_remain3_1393;
address_decode_4 decoder_3_1393 = address_decode_4(addr_selector2_87[1],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1393,addr_remain3_1393);


wire[15:0] addr_selector3_1394;
wire[15:0] addr_remain3_1394;
address_decode_4 decoder_3_1394 = address_decode_4(addr_selector2_87[2],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1394,addr_remain3_1394);


wire[15:0] addr_selector3_1395;
wire[15:0] addr_remain3_1395;
address_decode_4 decoder_3_1395 = address_decode_4(addr_selector2_87[3],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1395,addr_remain3_1395);


wire[15:0] addr_selector3_1396;
wire[15:0] addr_remain3_1396;
address_decode_4 decoder_3_1396 = address_decode_4(addr_selector2_87[4],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1396,addr_remain3_1396);


wire[15:0] addr_selector3_1397;
wire[15:0] addr_remain3_1397;
address_decode_4 decoder_3_1397 = address_decode_4(addr_selector2_87[5],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1397,addr_remain3_1397);


wire[15:0] addr_selector3_1398;
wire[15:0] addr_remain3_1398;
address_decode_4 decoder_3_1398 = address_decode_4(addr_selector2_87[6],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1398,addr_remain3_1398);


wire[15:0] addr_selector3_1399;
wire[15:0] addr_remain3_1399;
address_decode_4 decoder_3_1399 = address_decode_4(addr_selector2_87[7],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1399,addr_remain3_1399);


wire[15:0] addr_selector3_1400;
wire[15:0] addr_remain3_1400;
address_decode_4 decoder_3_1400 = address_decode_4(addr_selector2_87[8],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1400,addr_remain3_1400);


wire[15:0] addr_selector3_1401;
wire[15:0] addr_remain3_1401;
address_decode_4 decoder_3_1401 = address_decode_4(addr_selector2_87[9],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1401,addr_remain3_1401);


wire[15:0] addr_selector3_1402;
wire[15:0] addr_remain3_1402;
address_decode_4 decoder_3_1402 = address_decode_4(addr_selector2_87[10],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1402,addr_remain3_1402);


wire[15:0] addr_selector3_1403;
wire[15:0] addr_remain3_1403;
address_decode_4 decoder_3_1403 = address_decode_4(addr_selector2_87[11],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1403,addr_remain3_1403);


wire[15:0] addr_selector3_1404;
wire[15:0] addr_remain3_1404;
address_decode_4 decoder_3_1404 = address_decode_4(addr_selector2_87[12],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1404,addr_remain3_1404);


wire[15:0] addr_selector3_1405;
wire[15:0] addr_remain3_1405;
address_decode_4 decoder_3_1405 = address_decode_4(addr_selector2_87[13],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1405,addr_remain3_1405);


wire[15:0] addr_selector3_1406;
wire[15:0] addr_remain3_1406;
address_decode_4 decoder_3_1406 = address_decode_4(addr_selector2_87[14],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1406,addr_remain3_1406);


wire[15:0] addr_selector3_1407;
wire[15:0] addr_remain3_1407;
address_decode_4 decoder_3_1407 = address_decode_4(addr_selector2_87[15],addr_remain2_87[15:0],addr_remain2_87,addr_selector3_1407,addr_remain3_1407);


wire[15:0] addr_selector3_1408;
wire[15:0] addr_remain3_1408;
address_decode_4 decoder_3_1408 = address_decode_4(addr_selector2_88[0],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1408,addr_remain3_1408);


wire[15:0] addr_selector3_1409;
wire[15:0] addr_remain3_1409;
address_decode_4 decoder_3_1409 = address_decode_4(addr_selector2_88[1],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1409,addr_remain3_1409);


wire[15:0] addr_selector3_1410;
wire[15:0] addr_remain3_1410;
address_decode_4 decoder_3_1410 = address_decode_4(addr_selector2_88[2],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1410,addr_remain3_1410);


wire[15:0] addr_selector3_1411;
wire[15:0] addr_remain3_1411;
address_decode_4 decoder_3_1411 = address_decode_4(addr_selector2_88[3],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1411,addr_remain3_1411);


wire[15:0] addr_selector3_1412;
wire[15:0] addr_remain3_1412;
address_decode_4 decoder_3_1412 = address_decode_4(addr_selector2_88[4],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1412,addr_remain3_1412);


wire[15:0] addr_selector3_1413;
wire[15:0] addr_remain3_1413;
address_decode_4 decoder_3_1413 = address_decode_4(addr_selector2_88[5],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1413,addr_remain3_1413);


wire[15:0] addr_selector3_1414;
wire[15:0] addr_remain3_1414;
address_decode_4 decoder_3_1414 = address_decode_4(addr_selector2_88[6],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1414,addr_remain3_1414);


wire[15:0] addr_selector3_1415;
wire[15:0] addr_remain3_1415;
address_decode_4 decoder_3_1415 = address_decode_4(addr_selector2_88[7],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1415,addr_remain3_1415);


wire[15:0] addr_selector3_1416;
wire[15:0] addr_remain3_1416;
address_decode_4 decoder_3_1416 = address_decode_4(addr_selector2_88[8],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1416,addr_remain3_1416);


wire[15:0] addr_selector3_1417;
wire[15:0] addr_remain3_1417;
address_decode_4 decoder_3_1417 = address_decode_4(addr_selector2_88[9],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1417,addr_remain3_1417);


wire[15:0] addr_selector3_1418;
wire[15:0] addr_remain3_1418;
address_decode_4 decoder_3_1418 = address_decode_4(addr_selector2_88[10],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1418,addr_remain3_1418);


wire[15:0] addr_selector3_1419;
wire[15:0] addr_remain3_1419;
address_decode_4 decoder_3_1419 = address_decode_4(addr_selector2_88[11],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1419,addr_remain3_1419);


wire[15:0] addr_selector3_1420;
wire[15:0] addr_remain3_1420;
address_decode_4 decoder_3_1420 = address_decode_4(addr_selector2_88[12],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1420,addr_remain3_1420);


wire[15:0] addr_selector3_1421;
wire[15:0] addr_remain3_1421;
address_decode_4 decoder_3_1421 = address_decode_4(addr_selector2_88[13],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1421,addr_remain3_1421);


wire[15:0] addr_selector3_1422;
wire[15:0] addr_remain3_1422;
address_decode_4 decoder_3_1422 = address_decode_4(addr_selector2_88[14],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1422,addr_remain3_1422);


wire[15:0] addr_selector3_1423;
wire[15:0] addr_remain3_1423;
address_decode_4 decoder_3_1423 = address_decode_4(addr_selector2_88[15],addr_remain2_88[15:0],addr_remain2_88,addr_selector3_1423,addr_remain3_1423);


wire[15:0] addr_selector3_1424;
wire[15:0] addr_remain3_1424;
address_decode_4 decoder_3_1424 = address_decode_4(addr_selector2_89[0],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1424,addr_remain3_1424);


wire[15:0] addr_selector3_1425;
wire[15:0] addr_remain3_1425;
address_decode_4 decoder_3_1425 = address_decode_4(addr_selector2_89[1],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1425,addr_remain3_1425);


wire[15:0] addr_selector3_1426;
wire[15:0] addr_remain3_1426;
address_decode_4 decoder_3_1426 = address_decode_4(addr_selector2_89[2],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1426,addr_remain3_1426);


wire[15:0] addr_selector3_1427;
wire[15:0] addr_remain3_1427;
address_decode_4 decoder_3_1427 = address_decode_4(addr_selector2_89[3],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1427,addr_remain3_1427);


wire[15:0] addr_selector3_1428;
wire[15:0] addr_remain3_1428;
address_decode_4 decoder_3_1428 = address_decode_4(addr_selector2_89[4],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1428,addr_remain3_1428);


wire[15:0] addr_selector3_1429;
wire[15:0] addr_remain3_1429;
address_decode_4 decoder_3_1429 = address_decode_4(addr_selector2_89[5],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1429,addr_remain3_1429);


wire[15:0] addr_selector3_1430;
wire[15:0] addr_remain3_1430;
address_decode_4 decoder_3_1430 = address_decode_4(addr_selector2_89[6],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1430,addr_remain3_1430);


wire[15:0] addr_selector3_1431;
wire[15:0] addr_remain3_1431;
address_decode_4 decoder_3_1431 = address_decode_4(addr_selector2_89[7],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1431,addr_remain3_1431);


wire[15:0] addr_selector3_1432;
wire[15:0] addr_remain3_1432;
address_decode_4 decoder_3_1432 = address_decode_4(addr_selector2_89[8],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1432,addr_remain3_1432);


wire[15:0] addr_selector3_1433;
wire[15:0] addr_remain3_1433;
address_decode_4 decoder_3_1433 = address_decode_4(addr_selector2_89[9],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1433,addr_remain3_1433);


wire[15:0] addr_selector3_1434;
wire[15:0] addr_remain3_1434;
address_decode_4 decoder_3_1434 = address_decode_4(addr_selector2_89[10],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1434,addr_remain3_1434);


wire[15:0] addr_selector3_1435;
wire[15:0] addr_remain3_1435;
address_decode_4 decoder_3_1435 = address_decode_4(addr_selector2_89[11],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1435,addr_remain3_1435);


wire[15:0] addr_selector3_1436;
wire[15:0] addr_remain3_1436;
address_decode_4 decoder_3_1436 = address_decode_4(addr_selector2_89[12],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1436,addr_remain3_1436);


wire[15:0] addr_selector3_1437;
wire[15:0] addr_remain3_1437;
address_decode_4 decoder_3_1437 = address_decode_4(addr_selector2_89[13],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1437,addr_remain3_1437);


wire[15:0] addr_selector3_1438;
wire[15:0] addr_remain3_1438;
address_decode_4 decoder_3_1438 = address_decode_4(addr_selector2_89[14],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1438,addr_remain3_1438);


wire[15:0] addr_selector3_1439;
wire[15:0] addr_remain3_1439;
address_decode_4 decoder_3_1439 = address_decode_4(addr_selector2_89[15],addr_remain2_89[15:0],addr_remain2_89,addr_selector3_1439,addr_remain3_1439);


wire[15:0] addr_selector3_1440;
wire[15:0] addr_remain3_1440;
address_decode_4 decoder_3_1440 = address_decode_4(addr_selector2_90[0],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1440,addr_remain3_1440);


wire[15:0] addr_selector3_1441;
wire[15:0] addr_remain3_1441;
address_decode_4 decoder_3_1441 = address_decode_4(addr_selector2_90[1],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1441,addr_remain3_1441);


wire[15:0] addr_selector3_1442;
wire[15:0] addr_remain3_1442;
address_decode_4 decoder_3_1442 = address_decode_4(addr_selector2_90[2],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1442,addr_remain3_1442);


wire[15:0] addr_selector3_1443;
wire[15:0] addr_remain3_1443;
address_decode_4 decoder_3_1443 = address_decode_4(addr_selector2_90[3],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1443,addr_remain3_1443);


wire[15:0] addr_selector3_1444;
wire[15:0] addr_remain3_1444;
address_decode_4 decoder_3_1444 = address_decode_4(addr_selector2_90[4],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1444,addr_remain3_1444);


wire[15:0] addr_selector3_1445;
wire[15:0] addr_remain3_1445;
address_decode_4 decoder_3_1445 = address_decode_4(addr_selector2_90[5],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1445,addr_remain3_1445);


wire[15:0] addr_selector3_1446;
wire[15:0] addr_remain3_1446;
address_decode_4 decoder_3_1446 = address_decode_4(addr_selector2_90[6],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1446,addr_remain3_1446);


wire[15:0] addr_selector3_1447;
wire[15:0] addr_remain3_1447;
address_decode_4 decoder_3_1447 = address_decode_4(addr_selector2_90[7],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1447,addr_remain3_1447);


wire[15:0] addr_selector3_1448;
wire[15:0] addr_remain3_1448;
address_decode_4 decoder_3_1448 = address_decode_4(addr_selector2_90[8],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1448,addr_remain3_1448);


wire[15:0] addr_selector3_1449;
wire[15:0] addr_remain3_1449;
address_decode_4 decoder_3_1449 = address_decode_4(addr_selector2_90[9],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1449,addr_remain3_1449);


wire[15:0] addr_selector3_1450;
wire[15:0] addr_remain3_1450;
address_decode_4 decoder_3_1450 = address_decode_4(addr_selector2_90[10],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1450,addr_remain3_1450);


wire[15:0] addr_selector3_1451;
wire[15:0] addr_remain3_1451;
address_decode_4 decoder_3_1451 = address_decode_4(addr_selector2_90[11],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1451,addr_remain3_1451);


wire[15:0] addr_selector3_1452;
wire[15:0] addr_remain3_1452;
address_decode_4 decoder_3_1452 = address_decode_4(addr_selector2_90[12],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1452,addr_remain3_1452);


wire[15:0] addr_selector3_1453;
wire[15:0] addr_remain3_1453;
address_decode_4 decoder_3_1453 = address_decode_4(addr_selector2_90[13],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1453,addr_remain3_1453);


wire[15:0] addr_selector3_1454;
wire[15:0] addr_remain3_1454;
address_decode_4 decoder_3_1454 = address_decode_4(addr_selector2_90[14],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1454,addr_remain3_1454);


wire[15:0] addr_selector3_1455;
wire[15:0] addr_remain3_1455;
address_decode_4 decoder_3_1455 = address_decode_4(addr_selector2_90[15],addr_remain2_90[15:0],addr_remain2_90,addr_selector3_1455,addr_remain3_1455);


wire[15:0] addr_selector3_1456;
wire[15:0] addr_remain3_1456;
address_decode_4 decoder_3_1456 = address_decode_4(addr_selector2_91[0],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1456,addr_remain3_1456);


wire[15:0] addr_selector3_1457;
wire[15:0] addr_remain3_1457;
address_decode_4 decoder_3_1457 = address_decode_4(addr_selector2_91[1],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1457,addr_remain3_1457);


wire[15:0] addr_selector3_1458;
wire[15:0] addr_remain3_1458;
address_decode_4 decoder_3_1458 = address_decode_4(addr_selector2_91[2],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1458,addr_remain3_1458);


wire[15:0] addr_selector3_1459;
wire[15:0] addr_remain3_1459;
address_decode_4 decoder_3_1459 = address_decode_4(addr_selector2_91[3],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1459,addr_remain3_1459);


wire[15:0] addr_selector3_1460;
wire[15:0] addr_remain3_1460;
address_decode_4 decoder_3_1460 = address_decode_4(addr_selector2_91[4],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1460,addr_remain3_1460);


wire[15:0] addr_selector3_1461;
wire[15:0] addr_remain3_1461;
address_decode_4 decoder_3_1461 = address_decode_4(addr_selector2_91[5],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1461,addr_remain3_1461);


wire[15:0] addr_selector3_1462;
wire[15:0] addr_remain3_1462;
address_decode_4 decoder_3_1462 = address_decode_4(addr_selector2_91[6],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1462,addr_remain3_1462);


wire[15:0] addr_selector3_1463;
wire[15:0] addr_remain3_1463;
address_decode_4 decoder_3_1463 = address_decode_4(addr_selector2_91[7],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1463,addr_remain3_1463);


wire[15:0] addr_selector3_1464;
wire[15:0] addr_remain3_1464;
address_decode_4 decoder_3_1464 = address_decode_4(addr_selector2_91[8],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1464,addr_remain3_1464);


wire[15:0] addr_selector3_1465;
wire[15:0] addr_remain3_1465;
address_decode_4 decoder_3_1465 = address_decode_4(addr_selector2_91[9],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1465,addr_remain3_1465);


wire[15:0] addr_selector3_1466;
wire[15:0] addr_remain3_1466;
address_decode_4 decoder_3_1466 = address_decode_4(addr_selector2_91[10],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1466,addr_remain3_1466);


wire[15:0] addr_selector3_1467;
wire[15:0] addr_remain3_1467;
address_decode_4 decoder_3_1467 = address_decode_4(addr_selector2_91[11],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1467,addr_remain3_1467);


wire[15:0] addr_selector3_1468;
wire[15:0] addr_remain3_1468;
address_decode_4 decoder_3_1468 = address_decode_4(addr_selector2_91[12],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1468,addr_remain3_1468);


wire[15:0] addr_selector3_1469;
wire[15:0] addr_remain3_1469;
address_decode_4 decoder_3_1469 = address_decode_4(addr_selector2_91[13],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1469,addr_remain3_1469);


wire[15:0] addr_selector3_1470;
wire[15:0] addr_remain3_1470;
address_decode_4 decoder_3_1470 = address_decode_4(addr_selector2_91[14],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1470,addr_remain3_1470);


wire[15:0] addr_selector3_1471;
wire[15:0] addr_remain3_1471;
address_decode_4 decoder_3_1471 = address_decode_4(addr_selector2_91[15],addr_remain2_91[15:0],addr_remain2_91,addr_selector3_1471,addr_remain3_1471);


wire[15:0] addr_selector3_1472;
wire[15:0] addr_remain3_1472;
address_decode_4 decoder_3_1472 = address_decode_4(addr_selector2_92[0],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1472,addr_remain3_1472);


wire[15:0] addr_selector3_1473;
wire[15:0] addr_remain3_1473;
address_decode_4 decoder_3_1473 = address_decode_4(addr_selector2_92[1],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1473,addr_remain3_1473);


wire[15:0] addr_selector3_1474;
wire[15:0] addr_remain3_1474;
address_decode_4 decoder_3_1474 = address_decode_4(addr_selector2_92[2],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1474,addr_remain3_1474);


wire[15:0] addr_selector3_1475;
wire[15:0] addr_remain3_1475;
address_decode_4 decoder_3_1475 = address_decode_4(addr_selector2_92[3],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1475,addr_remain3_1475);


wire[15:0] addr_selector3_1476;
wire[15:0] addr_remain3_1476;
address_decode_4 decoder_3_1476 = address_decode_4(addr_selector2_92[4],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1476,addr_remain3_1476);


wire[15:0] addr_selector3_1477;
wire[15:0] addr_remain3_1477;
address_decode_4 decoder_3_1477 = address_decode_4(addr_selector2_92[5],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1477,addr_remain3_1477);


wire[15:0] addr_selector3_1478;
wire[15:0] addr_remain3_1478;
address_decode_4 decoder_3_1478 = address_decode_4(addr_selector2_92[6],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1478,addr_remain3_1478);


wire[15:0] addr_selector3_1479;
wire[15:0] addr_remain3_1479;
address_decode_4 decoder_3_1479 = address_decode_4(addr_selector2_92[7],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1479,addr_remain3_1479);


wire[15:0] addr_selector3_1480;
wire[15:0] addr_remain3_1480;
address_decode_4 decoder_3_1480 = address_decode_4(addr_selector2_92[8],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1480,addr_remain3_1480);


wire[15:0] addr_selector3_1481;
wire[15:0] addr_remain3_1481;
address_decode_4 decoder_3_1481 = address_decode_4(addr_selector2_92[9],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1481,addr_remain3_1481);


wire[15:0] addr_selector3_1482;
wire[15:0] addr_remain3_1482;
address_decode_4 decoder_3_1482 = address_decode_4(addr_selector2_92[10],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1482,addr_remain3_1482);


wire[15:0] addr_selector3_1483;
wire[15:0] addr_remain3_1483;
address_decode_4 decoder_3_1483 = address_decode_4(addr_selector2_92[11],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1483,addr_remain3_1483);


wire[15:0] addr_selector3_1484;
wire[15:0] addr_remain3_1484;
address_decode_4 decoder_3_1484 = address_decode_4(addr_selector2_92[12],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1484,addr_remain3_1484);


wire[15:0] addr_selector3_1485;
wire[15:0] addr_remain3_1485;
address_decode_4 decoder_3_1485 = address_decode_4(addr_selector2_92[13],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1485,addr_remain3_1485);


wire[15:0] addr_selector3_1486;
wire[15:0] addr_remain3_1486;
address_decode_4 decoder_3_1486 = address_decode_4(addr_selector2_92[14],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1486,addr_remain3_1486);


wire[15:0] addr_selector3_1487;
wire[15:0] addr_remain3_1487;
address_decode_4 decoder_3_1487 = address_decode_4(addr_selector2_92[15],addr_remain2_92[15:0],addr_remain2_92,addr_selector3_1487,addr_remain3_1487);


wire[15:0] addr_selector3_1488;
wire[15:0] addr_remain3_1488;
address_decode_4 decoder_3_1488 = address_decode_4(addr_selector2_93[0],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1488,addr_remain3_1488);


wire[15:0] addr_selector3_1489;
wire[15:0] addr_remain3_1489;
address_decode_4 decoder_3_1489 = address_decode_4(addr_selector2_93[1],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1489,addr_remain3_1489);


wire[15:0] addr_selector3_1490;
wire[15:0] addr_remain3_1490;
address_decode_4 decoder_3_1490 = address_decode_4(addr_selector2_93[2],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1490,addr_remain3_1490);


wire[15:0] addr_selector3_1491;
wire[15:0] addr_remain3_1491;
address_decode_4 decoder_3_1491 = address_decode_4(addr_selector2_93[3],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1491,addr_remain3_1491);


wire[15:0] addr_selector3_1492;
wire[15:0] addr_remain3_1492;
address_decode_4 decoder_3_1492 = address_decode_4(addr_selector2_93[4],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1492,addr_remain3_1492);


wire[15:0] addr_selector3_1493;
wire[15:0] addr_remain3_1493;
address_decode_4 decoder_3_1493 = address_decode_4(addr_selector2_93[5],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1493,addr_remain3_1493);


wire[15:0] addr_selector3_1494;
wire[15:0] addr_remain3_1494;
address_decode_4 decoder_3_1494 = address_decode_4(addr_selector2_93[6],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1494,addr_remain3_1494);


wire[15:0] addr_selector3_1495;
wire[15:0] addr_remain3_1495;
address_decode_4 decoder_3_1495 = address_decode_4(addr_selector2_93[7],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1495,addr_remain3_1495);


wire[15:0] addr_selector3_1496;
wire[15:0] addr_remain3_1496;
address_decode_4 decoder_3_1496 = address_decode_4(addr_selector2_93[8],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1496,addr_remain3_1496);


wire[15:0] addr_selector3_1497;
wire[15:0] addr_remain3_1497;
address_decode_4 decoder_3_1497 = address_decode_4(addr_selector2_93[9],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1497,addr_remain3_1497);


wire[15:0] addr_selector3_1498;
wire[15:0] addr_remain3_1498;
address_decode_4 decoder_3_1498 = address_decode_4(addr_selector2_93[10],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1498,addr_remain3_1498);


wire[15:0] addr_selector3_1499;
wire[15:0] addr_remain3_1499;
address_decode_4 decoder_3_1499 = address_decode_4(addr_selector2_93[11],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1499,addr_remain3_1499);


wire[15:0] addr_selector3_1500;
wire[15:0] addr_remain3_1500;
address_decode_4 decoder_3_1500 = address_decode_4(addr_selector2_93[12],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1500,addr_remain3_1500);


wire[15:0] addr_selector3_1501;
wire[15:0] addr_remain3_1501;
address_decode_4 decoder_3_1501 = address_decode_4(addr_selector2_93[13],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1501,addr_remain3_1501);


wire[15:0] addr_selector3_1502;
wire[15:0] addr_remain3_1502;
address_decode_4 decoder_3_1502 = address_decode_4(addr_selector2_93[14],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1502,addr_remain3_1502);


wire[15:0] addr_selector3_1503;
wire[15:0] addr_remain3_1503;
address_decode_4 decoder_3_1503 = address_decode_4(addr_selector2_93[15],addr_remain2_93[15:0],addr_remain2_93,addr_selector3_1503,addr_remain3_1503);


wire[15:0] addr_selector3_1504;
wire[15:0] addr_remain3_1504;
address_decode_4 decoder_3_1504 = address_decode_4(addr_selector2_94[0],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1504,addr_remain3_1504);


wire[15:0] addr_selector3_1505;
wire[15:0] addr_remain3_1505;
address_decode_4 decoder_3_1505 = address_decode_4(addr_selector2_94[1],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1505,addr_remain3_1505);


wire[15:0] addr_selector3_1506;
wire[15:0] addr_remain3_1506;
address_decode_4 decoder_3_1506 = address_decode_4(addr_selector2_94[2],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1506,addr_remain3_1506);


wire[15:0] addr_selector3_1507;
wire[15:0] addr_remain3_1507;
address_decode_4 decoder_3_1507 = address_decode_4(addr_selector2_94[3],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1507,addr_remain3_1507);


wire[15:0] addr_selector3_1508;
wire[15:0] addr_remain3_1508;
address_decode_4 decoder_3_1508 = address_decode_4(addr_selector2_94[4],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1508,addr_remain3_1508);


wire[15:0] addr_selector3_1509;
wire[15:0] addr_remain3_1509;
address_decode_4 decoder_3_1509 = address_decode_4(addr_selector2_94[5],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1509,addr_remain3_1509);


wire[15:0] addr_selector3_1510;
wire[15:0] addr_remain3_1510;
address_decode_4 decoder_3_1510 = address_decode_4(addr_selector2_94[6],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1510,addr_remain3_1510);


wire[15:0] addr_selector3_1511;
wire[15:0] addr_remain3_1511;
address_decode_4 decoder_3_1511 = address_decode_4(addr_selector2_94[7],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1511,addr_remain3_1511);


wire[15:0] addr_selector3_1512;
wire[15:0] addr_remain3_1512;
address_decode_4 decoder_3_1512 = address_decode_4(addr_selector2_94[8],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1512,addr_remain3_1512);


wire[15:0] addr_selector3_1513;
wire[15:0] addr_remain3_1513;
address_decode_4 decoder_3_1513 = address_decode_4(addr_selector2_94[9],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1513,addr_remain3_1513);


wire[15:0] addr_selector3_1514;
wire[15:0] addr_remain3_1514;
address_decode_4 decoder_3_1514 = address_decode_4(addr_selector2_94[10],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1514,addr_remain3_1514);


wire[15:0] addr_selector3_1515;
wire[15:0] addr_remain3_1515;
address_decode_4 decoder_3_1515 = address_decode_4(addr_selector2_94[11],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1515,addr_remain3_1515);


wire[15:0] addr_selector3_1516;
wire[15:0] addr_remain3_1516;
address_decode_4 decoder_3_1516 = address_decode_4(addr_selector2_94[12],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1516,addr_remain3_1516);


wire[15:0] addr_selector3_1517;
wire[15:0] addr_remain3_1517;
address_decode_4 decoder_3_1517 = address_decode_4(addr_selector2_94[13],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1517,addr_remain3_1517);


wire[15:0] addr_selector3_1518;
wire[15:0] addr_remain3_1518;
address_decode_4 decoder_3_1518 = address_decode_4(addr_selector2_94[14],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1518,addr_remain3_1518);


wire[15:0] addr_selector3_1519;
wire[15:0] addr_remain3_1519;
address_decode_4 decoder_3_1519 = address_decode_4(addr_selector2_94[15],addr_remain2_94[15:0],addr_remain2_94,addr_selector3_1519,addr_remain3_1519);


wire[15:0] addr_selector3_1520;
wire[15:0] addr_remain3_1520;
address_decode_4 decoder_3_1520 = address_decode_4(addr_selector2_95[0],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1520,addr_remain3_1520);


wire[15:0] addr_selector3_1521;
wire[15:0] addr_remain3_1521;
address_decode_4 decoder_3_1521 = address_decode_4(addr_selector2_95[1],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1521,addr_remain3_1521);


wire[15:0] addr_selector3_1522;
wire[15:0] addr_remain3_1522;
address_decode_4 decoder_3_1522 = address_decode_4(addr_selector2_95[2],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1522,addr_remain3_1522);


wire[15:0] addr_selector3_1523;
wire[15:0] addr_remain3_1523;
address_decode_4 decoder_3_1523 = address_decode_4(addr_selector2_95[3],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1523,addr_remain3_1523);


wire[15:0] addr_selector3_1524;
wire[15:0] addr_remain3_1524;
address_decode_4 decoder_3_1524 = address_decode_4(addr_selector2_95[4],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1524,addr_remain3_1524);


wire[15:0] addr_selector3_1525;
wire[15:0] addr_remain3_1525;
address_decode_4 decoder_3_1525 = address_decode_4(addr_selector2_95[5],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1525,addr_remain3_1525);


wire[15:0] addr_selector3_1526;
wire[15:0] addr_remain3_1526;
address_decode_4 decoder_3_1526 = address_decode_4(addr_selector2_95[6],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1526,addr_remain3_1526);


wire[15:0] addr_selector3_1527;
wire[15:0] addr_remain3_1527;
address_decode_4 decoder_3_1527 = address_decode_4(addr_selector2_95[7],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1527,addr_remain3_1527);


wire[15:0] addr_selector3_1528;
wire[15:0] addr_remain3_1528;
address_decode_4 decoder_3_1528 = address_decode_4(addr_selector2_95[8],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1528,addr_remain3_1528);


wire[15:0] addr_selector3_1529;
wire[15:0] addr_remain3_1529;
address_decode_4 decoder_3_1529 = address_decode_4(addr_selector2_95[9],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1529,addr_remain3_1529);


wire[15:0] addr_selector3_1530;
wire[15:0] addr_remain3_1530;
address_decode_4 decoder_3_1530 = address_decode_4(addr_selector2_95[10],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1530,addr_remain3_1530);


wire[15:0] addr_selector3_1531;
wire[15:0] addr_remain3_1531;
address_decode_4 decoder_3_1531 = address_decode_4(addr_selector2_95[11],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1531,addr_remain3_1531);


wire[15:0] addr_selector3_1532;
wire[15:0] addr_remain3_1532;
address_decode_4 decoder_3_1532 = address_decode_4(addr_selector2_95[12],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1532,addr_remain3_1532);


wire[15:0] addr_selector3_1533;
wire[15:0] addr_remain3_1533;
address_decode_4 decoder_3_1533 = address_decode_4(addr_selector2_95[13],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1533,addr_remain3_1533);


wire[15:0] addr_selector3_1534;
wire[15:0] addr_remain3_1534;
address_decode_4 decoder_3_1534 = address_decode_4(addr_selector2_95[14],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1534,addr_remain3_1534);


wire[15:0] addr_selector3_1535;
wire[15:0] addr_remain3_1535;
address_decode_4 decoder_3_1535 = address_decode_4(addr_selector2_95[15],addr_remain2_95[15:0],addr_remain2_95,addr_selector3_1535,addr_remain3_1535);


wire[15:0] addr_selector3_1536;
wire[15:0] addr_remain3_1536;
address_decode_4 decoder_3_1536 = address_decode_4(addr_selector2_96[0],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1536,addr_remain3_1536);


wire[15:0] addr_selector3_1537;
wire[15:0] addr_remain3_1537;
address_decode_4 decoder_3_1537 = address_decode_4(addr_selector2_96[1],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1537,addr_remain3_1537);


wire[15:0] addr_selector3_1538;
wire[15:0] addr_remain3_1538;
address_decode_4 decoder_3_1538 = address_decode_4(addr_selector2_96[2],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1538,addr_remain3_1538);


wire[15:0] addr_selector3_1539;
wire[15:0] addr_remain3_1539;
address_decode_4 decoder_3_1539 = address_decode_4(addr_selector2_96[3],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1539,addr_remain3_1539);


wire[15:0] addr_selector3_1540;
wire[15:0] addr_remain3_1540;
address_decode_4 decoder_3_1540 = address_decode_4(addr_selector2_96[4],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1540,addr_remain3_1540);


wire[15:0] addr_selector3_1541;
wire[15:0] addr_remain3_1541;
address_decode_4 decoder_3_1541 = address_decode_4(addr_selector2_96[5],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1541,addr_remain3_1541);


wire[15:0] addr_selector3_1542;
wire[15:0] addr_remain3_1542;
address_decode_4 decoder_3_1542 = address_decode_4(addr_selector2_96[6],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1542,addr_remain3_1542);


wire[15:0] addr_selector3_1543;
wire[15:0] addr_remain3_1543;
address_decode_4 decoder_3_1543 = address_decode_4(addr_selector2_96[7],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1543,addr_remain3_1543);


wire[15:0] addr_selector3_1544;
wire[15:0] addr_remain3_1544;
address_decode_4 decoder_3_1544 = address_decode_4(addr_selector2_96[8],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1544,addr_remain3_1544);


wire[15:0] addr_selector3_1545;
wire[15:0] addr_remain3_1545;
address_decode_4 decoder_3_1545 = address_decode_4(addr_selector2_96[9],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1545,addr_remain3_1545);


wire[15:0] addr_selector3_1546;
wire[15:0] addr_remain3_1546;
address_decode_4 decoder_3_1546 = address_decode_4(addr_selector2_96[10],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1546,addr_remain3_1546);


wire[15:0] addr_selector3_1547;
wire[15:0] addr_remain3_1547;
address_decode_4 decoder_3_1547 = address_decode_4(addr_selector2_96[11],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1547,addr_remain3_1547);


wire[15:0] addr_selector3_1548;
wire[15:0] addr_remain3_1548;
address_decode_4 decoder_3_1548 = address_decode_4(addr_selector2_96[12],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1548,addr_remain3_1548);


wire[15:0] addr_selector3_1549;
wire[15:0] addr_remain3_1549;
address_decode_4 decoder_3_1549 = address_decode_4(addr_selector2_96[13],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1549,addr_remain3_1549);


wire[15:0] addr_selector3_1550;
wire[15:0] addr_remain3_1550;
address_decode_4 decoder_3_1550 = address_decode_4(addr_selector2_96[14],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1550,addr_remain3_1550);


wire[15:0] addr_selector3_1551;
wire[15:0] addr_remain3_1551;
address_decode_4 decoder_3_1551 = address_decode_4(addr_selector2_96[15],addr_remain2_96[15:0],addr_remain2_96,addr_selector3_1551,addr_remain3_1551);


wire[15:0] addr_selector3_1552;
wire[15:0] addr_remain3_1552;
address_decode_4 decoder_3_1552 = address_decode_4(addr_selector2_97[0],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1552,addr_remain3_1552);


wire[15:0] addr_selector3_1553;
wire[15:0] addr_remain3_1553;
address_decode_4 decoder_3_1553 = address_decode_4(addr_selector2_97[1],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1553,addr_remain3_1553);


wire[15:0] addr_selector3_1554;
wire[15:0] addr_remain3_1554;
address_decode_4 decoder_3_1554 = address_decode_4(addr_selector2_97[2],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1554,addr_remain3_1554);


wire[15:0] addr_selector3_1555;
wire[15:0] addr_remain3_1555;
address_decode_4 decoder_3_1555 = address_decode_4(addr_selector2_97[3],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1555,addr_remain3_1555);


wire[15:0] addr_selector3_1556;
wire[15:0] addr_remain3_1556;
address_decode_4 decoder_3_1556 = address_decode_4(addr_selector2_97[4],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1556,addr_remain3_1556);


wire[15:0] addr_selector3_1557;
wire[15:0] addr_remain3_1557;
address_decode_4 decoder_3_1557 = address_decode_4(addr_selector2_97[5],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1557,addr_remain3_1557);


wire[15:0] addr_selector3_1558;
wire[15:0] addr_remain3_1558;
address_decode_4 decoder_3_1558 = address_decode_4(addr_selector2_97[6],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1558,addr_remain3_1558);


wire[15:0] addr_selector3_1559;
wire[15:0] addr_remain3_1559;
address_decode_4 decoder_3_1559 = address_decode_4(addr_selector2_97[7],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1559,addr_remain3_1559);


wire[15:0] addr_selector3_1560;
wire[15:0] addr_remain3_1560;
address_decode_4 decoder_3_1560 = address_decode_4(addr_selector2_97[8],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1560,addr_remain3_1560);


wire[15:0] addr_selector3_1561;
wire[15:0] addr_remain3_1561;
address_decode_4 decoder_3_1561 = address_decode_4(addr_selector2_97[9],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1561,addr_remain3_1561);


wire[15:0] addr_selector3_1562;
wire[15:0] addr_remain3_1562;
address_decode_4 decoder_3_1562 = address_decode_4(addr_selector2_97[10],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1562,addr_remain3_1562);


wire[15:0] addr_selector3_1563;
wire[15:0] addr_remain3_1563;
address_decode_4 decoder_3_1563 = address_decode_4(addr_selector2_97[11],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1563,addr_remain3_1563);


wire[15:0] addr_selector3_1564;
wire[15:0] addr_remain3_1564;
address_decode_4 decoder_3_1564 = address_decode_4(addr_selector2_97[12],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1564,addr_remain3_1564);


wire[15:0] addr_selector3_1565;
wire[15:0] addr_remain3_1565;
address_decode_4 decoder_3_1565 = address_decode_4(addr_selector2_97[13],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1565,addr_remain3_1565);


wire[15:0] addr_selector3_1566;
wire[15:0] addr_remain3_1566;
address_decode_4 decoder_3_1566 = address_decode_4(addr_selector2_97[14],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1566,addr_remain3_1566);


wire[15:0] addr_selector3_1567;
wire[15:0] addr_remain3_1567;
address_decode_4 decoder_3_1567 = address_decode_4(addr_selector2_97[15],addr_remain2_97[15:0],addr_remain2_97,addr_selector3_1567,addr_remain3_1567);


wire[15:0] addr_selector3_1568;
wire[15:0] addr_remain3_1568;
address_decode_4 decoder_3_1568 = address_decode_4(addr_selector2_98[0],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1568,addr_remain3_1568);


wire[15:0] addr_selector3_1569;
wire[15:0] addr_remain3_1569;
address_decode_4 decoder_3_1569 = address_decode_4(addr_selector2_98[1],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1569,addr_remain3_1569);


wire[15:0] addr_selector3_1570;
wire[15:0] addr_remain3_1570;
address_decode_4 decoder_3_1570 = address_decode_4(addr_selector2_98[2],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1570,addr_remain3_1570);


wire[15:0] addr_selector3_1571;
wire[15:0] addr_remain3_1571;
address_decode_4 decoder_3_1571 = address_decode_4(addr_selector2_98[3],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1571,addr_remain3_1571);


wire[15:0] addr_selector3_1572;
wire[15:0] addr_remain3_1572;
address_decode_4 decoder_3_1572 = address_decode_4(addr_selector2_98[4],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1572,addr_remain3_1572);


wire[15:0] addr_selector3_1573;
wire[15:0] addr_remain3_1573;
address_decode_4 decoder_3_1573 = address_decode_4(addr_selector2_98[5],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1573,addr_remain3_1573);


wire[15:0] addr_selector3_1574;
wire[15:0] addr_remain3_1574;
address_decode_4 decoder_3_1574 = address_decode_4(addr_selector2_98[6],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1574,addr_remain3_1574);


wire[15:0] addr_selector3_1575;
wire[15:0] addr_remain3_1575;
address_decode_4 decoder_3_1575 = address_decode_4(addr_selector2_98[7],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1575,addr_remain3_1575);


wire[15:0] addr_selector3_1576;
wire[15:0] addr_remain3_1576;
address_decode_4 decoder_3_1576 = address_decode_4(addr_selector2_98[8],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1576,addr_remain3_1576);


wire[15:0] addr_selector3_1577;
wire[15:0] addr_remain3_1577;
address_decode_4 decoder_3_1577 = address_decode_4(addr_selector2_98[9],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1577,addr_remain3_1577);


wire[15:0] addr_selector3_1578;
wire[15:0] addr_remain3_1578;
address_decode_4 decoder_3_1578 = address_decode_4(addr_selector2_98[10],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1578,addr_remain3_1578);


wire[15:0] addr_selector3_1579;
wire[15:0] addr_remain3_1579;
address_decode_4 decoder_3_1579 = address_decode_4(addr_selector2_98[11],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1579,addr_remain3_1579);


wire[15:0] addr_selector3_1580;
wire[15:0] addr_remain3_1580;
address_decode_4 decoder_3_1580 = address_decode_4(addr_selector2_98[12],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1580,addr_remain3_1580);


wire[15:0] addr_selector3_1581;
wire[15:0] addr_remain3_1581;
address_decode_4 decoder_3_1581 = address_decode_4(addr_selector2_98[13],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1581,addr_remain3_1581);


wire[15:0] addr_selector3_1582;
wire[15:0] addr_remain3_1582;
address_decode_4 decoder_3_1582 = address_decode_4(addr_selector2_98[14],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1582,addr_remain3_1582);


wire[15:0] addr_selector3_1583;
wire[15:0] addr_remain3_1583;
address_decode_4 decoder_3_1583 = address_decode_4(addr_selector2_98[15],addr_remain2_98[15:0],addr_remain2_98,addr_selector3_1583,addr_remain3_1583);


wire[15:0] addr_selector3_1584;
wire[15:0] addr_remain3_1584;
address_decode_4 decoder_3_1584 = address_decode_4(addr_selector2_99[0],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1584,addr_remain3_1584);


wire[15:0] addr_selector3_1585;
wire[15:0] addr_remain3_1585;
address_decode_4 decoder_3_1585 = address_decode_4(addr_selector2_99[1],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1585,addr_remain3_1585);


wire[15:0] addr_selector3_1586;
wire[15:0] addr_remain3_1586;
address_decode_4 decoder_3_1586 = address_decode_4(addr_selector2_99[2],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1586,addr_remain3_1586);


wire[15:0] addr_selector3_1587;
wire[15:0] addr_remain3_1587;
address_decode_4 decoder_3_1587 = address_decode_4(addr_selector2_99[3],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1587,addr_remain3_1587);


wire[15:0] addr_selector3_1588;
wire[15:0] addr_remain3_1588;
address_decode_4 decoder_3_1588 = address_decode_4(addr_selector2_99[4],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1588,addr_remain3_1588);


wire[15:0] addr_selector3_1589;
wire[15:0] addr_remain3_1589;
address_decode_4 decoder_3_1589 = address_decode_4(addr_selector2_99[5],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1589,addr_remain3_1589);


wire[15:0] addr_selector3_1590;
wire[15:0] addr_remain3_1590;
address_decode_4 decoder_3_1590 = address_decode_4(addr_selector2_99[6],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1590,addr_remain3_1590);


wire[15:0] addr_selector3_1591;
wire[15:0] addr_remain3_1591;
address_decode_4 decoder_3_1591 = address_decode_4(addr_selector2_99[7],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1591,addr_remain3_1591);


wire[15:0] addr_selector3_1592;
wire[15:0] addr_remain3_1592;
address_decode_4 decoder_3_1592 = address_decode_4(addr_selector2_99[8],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1592,addr_remain3_1592);


wire[15:0] addr_selector3_1593;
wire[15:0] addr_remain3_1593;
address_decode_4 decoder_3_1593 = address_decode_4(addr_selector2_99[9],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1593,addr_remain3_1593);


wire[15:0] addr_selector3_1594;
wire[15:0] addr_remain3_1594;
address_decode_4 decoder_3_1594 = address_decode_4(addr_selector2_99[10],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1594,addr_remain3_1594);


wire[15:0] addr_selector3_1595;
wire[15:0] addr_remain3_1595;
address_decode_4 decoder_3_1595 = address_decode_4(addr_selector2_99[11],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1595,addr_remain3_1595);


wire[15:0] addr_selector3_1596;
wire[15:0] addr_remain3_1596;
address_decode_4 decoder_3_1596 = address_decode_4(addr_selector2_99[12],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1596,addr_remain3_1596);


wire[15:0] addr_selector3_1597;
wire[15:0] addr_remain3_1597;
address_decode_4 decoder_3_1597 = address_decode_4(addr_selector2_99[13],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1597,addr_remain3_1597);


wire[15:0] addr_selector3_1598;
wire[15:0] addr_remain3_1598;
address_decode_4 decoder_3_1598 = address_decode_4(addr_selector2_99[14],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1598,addr_remain3_1598);


wire[15:0] addr_selector3_1599;
wire[15:0] addr_remain3_1599;
address_decode_4 decoder_3_1599 = address_decode_4(addr_selector2_99[15],addr_remain2_99[15:0],addr_remain2_99,addr_selector3_1599,addr_remain3_1599);


wire[15:0] addr_selector3_1600;
wire[15:0] addr_remain3_1600;
address_decode_4 decoder_3_1600 = address_decode_4(addr_selector2_100[0],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1600,addr_remain3_1600);


wire[15:0] addr_selector3_1601;
wire[15:0] addr_remain3_1601;
address_decode_4 decoder_3_1601 = address_decode_4(addr_selector2_100[1],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1601,addr_remain3_1601);


wire[15:0] addr_selector3_1602;
wire[15:0] addr_remain3_1602;
address_decode_4 decoder_3_1602 = address_decode_4(addr_selector2_100[2],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1602,addr_remain3_1602);


wire[15:0] addr_selector3_1603;
wire[15:0] addr_remain3_1603;
address_decode_4 decoder_3_1603 = address_decode_4(addr_selector2_100[3],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1603,addr_remain3_1603);


wire[15:0] addr_selector3_1604;
wire[15:0] addr_remain3_1604;
address_decode_4 decoder_3_1604 = address_decode_4(addr_selector2_100[4],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1604,addr_remain3_1604);


wire[15:0] addr_selector3_1605;
wire[15:0] addr_remain3_1605;
address_decode_4 decoder_3_1605 = address_decode_4(addr_selector2_100[5],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1605,addr_remain3_1605);


wire[15:0] addr_selector3_1606;
wire[15:0] addr_remain3_1606;
address_decode_4 decoder_3_1606 = address_decode_4(addr_selector2_100[6],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1606,addr_remain3_1606);


wire[15:0] addr_selector3_1607;
wire[15:0] addr_remain3_1607;
address_decode_4 decoder_3_1607 = address_decode_4(addr_selector2_100[7],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1607,addr_remain3_1607);


wire[15:0] addr_selector3_1608;
wire[15:0] addr_remain3_1608;
address_decode_4 decoder_3_1608 = address_decode_4(addr_selector2_100[8],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1608,addr_remain3_1608);


wire[15:0] addr_selector3_1609;
wire[15:0] addr_remain3_1609;
address_decode_4 decoder_3_1609 = address_decode_4(addr_selector2_100[9],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1609,addr_remain3_1609);


wire[15:0] addr_selector3_1610;
wire[15:0] addr_remain3_1610;
address_decode_4 decoder_3_1610 = address_decode_4(addr_selector2_100[10],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1610,addr_remain3_1610);


wire[15:0] addr_selector3_1611;
wire[15:0] addr_remain3_1611;
address_decode_4 decoder_3_1611 = address_decode_4(addr_selector2_100[11],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1611,addr_remain3_1611);


wire[15:0] addr_selector3_1612;
wire[15:0] addr_remain3_1612;
address_decode_4 decoder_3_1612 = address_decode_4(addr_selector2_100[12],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1612,addr_remain3_1612);


wire[15:0] addr_selector3_1613;
wire[15:0] addr_remain3_1613;
address_decode_4 decoder_3_1613 = address_decode_4(addr_selector2_100[13],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1613,addr_remain3_1613);


wire[15:0] addr_selector3_1614;
wire[15:0] addr_remain3_1614;
address_decode_4 decoder_3_1614 = address_decode_4(addr_selector2_100[14],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1614,addr_remain3_1614);


wire[15:0] addr_selector3_1615;
wire[15:0] addr_remain3_1615;
address_decode_4 decoder_3_1615 = address_decode_4(addr_selector2_100[15],addr_remain2_100[15:0],addr_remain2_100,addr_selector3_1615,addr_remain3_1615);


wire[15:0] addr_selector3_1616;
wire[15:0] addr_remain3_1616;
address_decode_4 decoder_3_1616 = address_decode_4(addr_selector2_101[0],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1616,addr_remain3_1616);


wire[15:0] addr_selector3_1617;
wire[15:0] addr_remain3_1617;
address_decode_4 decoder_3_1617 = address_decode_4(addr_selector2_101[1],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1617,addr_remain3_1617);


wire[15:0] addr_selector3_1618;
wire[15:0] addr_remain3_1618;
address_decode_4 decoder_3_1618 = address_decode_4(addr_selector2_101[2],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1618,addr_remain3_1618);


wire[15:0] addr_selector3_1619;
wire[15:0] addr_remain3_1619;
address_decode_4 decoder_3_1619 = address_decode_4(addr_selector2_101[3],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1619,addr_remain3_1619);


wire[15:0] addr_selector3_1620;
wire[15:0] addr_remain3_1620;
address_decode_4 decoder_3_1620 = address_decode_4(addr_selector2_101[4],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1620,addr_remain3_1620);


wire[15:0] addr_selector3_1621;
wire[15:0] addr_remain3_1621;
address_decode_4 decoder_3_1621 = address_decode_4(addr_selector2_101[5],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1621,addr_remain3_1621);


wire[15:0] addr_selector3_1622;
wire[15:0] addr_remain3_1622;
address_decode_4 decoder_3_1622 = address_decode_4(addr_selector2_101[6],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1622,addr_remain3_1622);


wire[15:0] addr_selector3_1623;
wire[15:0] addr_remain3_1623;
address_decode_4 decoder_3_1623 = address_decode_4(addr_selector2_101[7],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1623,addr_remain3_1623);


wire[15:0] addr_selector3_1624;
wire[15:0] addr_remain3_1624;
address_decode_4 decoder_3_1624 = address_decode_4(addr_selector2_101[8],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1624,addr_remain3_1624);


wire[15:0] addr_selector3_1625;
wire[15:0] addr_remain3_1625;
address_decode_4 decoder_3_1625 = address_decode_4(addr_selector2_101[9],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1625,addr_remain3_1625);


wire[15:0] addr_selector3_1626;
wire[15:0] addr_remain3_1626;
address_decode_4 decoder_3_1626 = address_decode_4(addr_selector2_101[10],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1626,addr_remain3_1626);


wire[15:0] addr_selector3_1627;
wire[15:0] addr_remain3_1627;
address_decode_4 decoder_3_1627 = address_decode_4(addr_selector2_101[11],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1627,addr_remain3_1627);


wire[15:0] addr_selector3_1628;
wire[15:0] addr_remain3_1628;
address_decode_4 decoder_3_1628 = address_decode_4(addr_selector2_101[12],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1628,addr_remain3_1628);


wire[15:0] addr_selector3_1629;
wire[15:0] addr_remain3_1629;
address_decode_4 decoder_3_1629 = address_decode_4(addr_selector2_101[13],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1629,addr_remain3_1629);


wire[15:0] addr_selector3_1630;
wire[15:0] addr_remain3_1630;
address_decode_4 decoder_3_1630 = address_decode_4(addr_selector2_101[14],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1630,addr_remain3_1630);


wire[15:0] addr_selector3_1631;
wire[15:0] addr_remain3_1631;
address_decode_4 decoder_3_1631 = address_decode_4(addr_selector2_101[15],addr_remain2_101[15:0],addr_remain2_101,addr_selector3_1631,addr_remain3_1631);


wire[15:0] addr_selector3_1632;
wire[15:0] addr_remain3_1632;
address_decode_4 decoder_3_1632 = address_decode_4(addr_selector2_102[0],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1632,addr_remain3_1632);


wire[15:0] addr_selector3_1633;
wire[15:0] addr_remain3_1633;
address_decode_4 decoder_3_1633 = address_decode_4(addr_selector2_102[1],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1633,addr_remain3_1633);


wire[15:0] addr_selector3_1634;
wire[15:0] addr_remain3_1634;
address_decode_4 decoder_3_1634 = address_decode_4(addr_selector2_102[2],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1634,addr_remain3_1634);


wire[15:0] addr_selector3_1635;
wire[15:0] addr_remain3_1635;
address_decode_4 decoder_3_1635 = address_decode_4(addr_selector2_102[3],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1635,addr_remain3_1635);


wire[15:0] addr_selector3_1636;
wire[15:0] addr_remain3_1636;
address_decode_4 decoder_3_1636 = address_decode_4(addr_selector2_102[4],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1636,addr_remain3_1636);


wire[15:0] addr_selector3_1637;
wire[15:0] addr_remain3_1637;
address_decode_4 decoder_3_1637 = address_decode_4(addr_selector2_102[5],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1637,addr_remain3_1637);


wire[15:0] addr_selector3_1638;
wire[15:0] addr_remain3_1638;
address_decode_4 decoder_3_1638 = address_decode_4(addr_selector2_102[6],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1638,addr_remain3_1638);


wire[15:0] addr_selector3_1639;
wire[15:0] addr_remain3_1639;
address_decode_4 decoder_3_1639 = address_decode_4(addr_selector2_102[7],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1639,addr_remain3_1639);


wire[15:0] addr_selector3_1640;
wire[15:0] addr_remain3_1640;
address_decode_4 decoder_3_1640 = address_decode_4(addr_selector2_102[8],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1640,addr_remain3_1640);


wire[15:0] addr_selector3_1641;
wire[15:0] addr_remain3_1641;
address_decode_4 decoder_3_1641 = address_decode_4(addr_selector2_102[9],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1641,addr_remain3_1641);


wire[15:0] addr_selector3_1642;
wire[15:0] addr_remain3_1642;
address_decode_4 decoder_3_1642 = address_decode_4(addr_selector2_102[10],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1642,addr_remain3_1642);


wire[15:0] addr_selector3_1643;
wire[15:0] addr_remain3_1643;
address_decode_4 decoder_3_1643 = address_decode_4(addr_selector2_102[11],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1643,addr_remain3_1643);


wire[15:0] addr_selector3_1644;
wire[15:0] addr_remain3_1644;
address_decode_4 decoder_3_1644 = address_decode_4(addr_selector2_102[12],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1644,addr_remain3_1644);


wire[15:0] addr_selector3_1645;
wire[15:0] addr_remain3_1645;
address_decode_4 decoder_3_1645 = address_decode_4(addr_selector2_102[13],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1645,addr_remain3_1645);


wire[15:0] addr_selector3_1646;
wire[15:0] addr_remain3_1646;
address_decode_4 decoder_3_1646 = address_decode_4(addr_selector2_102[14],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1646,addr_remain3_1646);


wire[15:0] addr_selector3_1647;
wire[15:0] addr_remain3_1647;
address_decode_4 decoder_3_1647 = address_decode_4(addr_selector2_102[15],addr_remain2_102[15:0],addr_remain2_102,addr_selector3_1647,addr_remain3_1647);


wire[15:0] addr_selector3_1648;
wire[15:0] addr_remain3_1648;
address_decode_4 decoder_3_1648 = address_decode_4(addr_selector2_103[0],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1648,addr_remain3_1648);


wire[15:0] addr_selector3_1649;
wire[15:0] addr_remain3_1649;
address_decode_4 decoder_3_1649 = address_decode_4(addr_selector2_103[1],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1649,addr_remain3_1649);


wire[15:0] addr_selector3_1650;
wire[15:0] addr_remain3_1650;
address_decode_4 decoder_3_1650 = address_decode_4(addr_selector2_103[2],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1650,addr_remain3_1650);


wire[15:0] addr_selector3_1651;
wire[15:0] addr_remain3_1651;
address_decode_4 decoder_3_1651 = address_decode_4(addr_selector2_103[3],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1651,addr_remain3_1651);


wire[15:0] addr_selector3_1652;
wire[15:0] addr_remain3_1652;
address_decode_4 decoder_3_1652 = address_decode_4(addr_selector2_103[4],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1652,addr_remain3_1652);


wire[15:0] addr_selector3_1653;
wire[15:0] addr_remain3_1653;
address_decode_4 decoder_3_1653 = address_decode_4(addr_selector2_103[5],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1653,addr_remain3_1653);


wire[15:0] addr_selector3_1654;
wire[15:0] addr_remain3_1654;
address_decode_4 decoder_3_1654 = address_decode_4(addr_selector2_103[6],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1654,addr_remain3_1654);


wire[15:0] addr_selector3_1655;
wire[15:0] addr_remain3_1655;
address_decode_4 decoder_3_1655 = address_decode_4(addr_selector2_103[7],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1655,addr_remain3_1655);


wire[15:0] addr_selector3_1656;
wire[15:0] addr_remain3_1656;
address_decode_4 decoder_3_1656 = address_decode_4(addr_selector2_103[8],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1656,addr_remain3_1656);


wire[15:0] addr_selector3_1657;
wire[15:0] addr_remain3_1657;
address_decode_4 decoder_3_1657 = address_decode_4(addr_selector2_103[9],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1657,addr_remain3_1657);


wire[15:0] addr_selector3_1658;
wire[15:0] addr_remain3_1658;
address_decode_4 decoder_3_1658 = address_decode_4(addr_selector2_103[10],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1658,addr_remain3_1658);


wire[15:0] addr_selector3_1659;
wire[15:0] addr_remain3_1659;
address_decode_4 decoder_3_1659 = address_decode_4(addr_selector2_103[11],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1659,addr_remain3_1659);


wire[15:0] addr_selector3_1660;
wire[15:0] addr_remain3_1660;
address_decode_4 decoder_3_1660 = address_decode_4(addr_selector2_103[12],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1660,addr_remain3_1660);


wire[15:0] addr_selector3_1661;
wire[15:0] addr_remain3_1661;
address_decode_4 decoder_3_1661 = address_decode_4(addr_selector2_103[13],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1661,addr_remain3_1661);


wire[15:0] addr_selector3_1662;
wire[15:0] addr_remain3_1662;
address_decode_4 decoder_3_1662 = address_decode_4(addr_selector2_103[14],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1662,addr_remain3_1662);


wire[15:0] addr_selector3_1663;
wire[15:0] addr_remain3_1663;
address_decode_4 decoder_3_1663 = address_decode_4(addr_selector2_103[15],addr_remain2_103[15:0],addr_remain2_103,addr_selector3_1663,addr_remain3_1663);


wire[15:0] addr_selector3_1664;
wire[15:0] addr_remain3_1664;
address_decode_4 decoder_3_1664 = address_decode_4(addr_selector2_104[0],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1664,addr_remain3_1664);


wire[15:0] addr_selector3_1665;
wire[15:0] addr_remain3_1665;
address_decode_4 decoder_3_1665 = address_decode_4(addr_selector2_104[1],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1665,addr_remain3_1665);


wire[15:0] addr_selector3_1666;
wire[15:0] addr_remain3_1666;
address_decode_4 decoder_3_1666 = address_decode_4(addr_selector2_104[2],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1666,addr_remain3_1666);


wire[15:0] addr_selector3_1667;
wire[15:0] addr_remain3_1667;
address_decode_4 decoder_3_1667 = address_decode_4(addr_selector2_104[3],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1667,addr_remain3_1667);


wire[15:0] addr_selector3_1668;
wire[15:0] addr_remain3_1668;
address_decode_4 decoder_3_1668 = address_decode_4(addr_selector2_104[4],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1668,addr_remain3_1668);


wire[15:0] addr_selector3_1669;
wire[15:0] addr_remain3_1669;
address_decode_4 decoder_3_1669 = address_decode_4(addr_selector2_104[5],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1669,addr_remain3_1669);


wire[15:0] addr_selector3_1670;
wire[15:0] addr_remain3_1670;
address_decode_4 decoder_3_1670 = address_decode_4(addr_selector2_104[6],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1670,addr_remain3_1670);


wire[15:0] addr_selector3_1671;
wire[15:0] addr_remain3_1671;
address_decode_4 decoder_3_1671 = address_decode_4(addr_selector2_104[7],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1671,addr_remain3_1671);


wire[15:0] addr_selector3_1672;
wire[15:0] addr_remain3_1672;
address_decode_4 decoder_3_1672 = address_decode_4(addr_selector2_104[8],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1672,addr_remain3_1672);


wire[15:0] addr_selector3_1673;
wire[15:0] addr_remain3_1673;
address_decode_4 decoder_3_1673 = address_decode_4(addr_selector2_104[9],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1673,addr_remain3_1673);


wire[15:0] addr_selector3_1674;
wire[15:0] addr_remain3_1674;
address_decode_4 decoder_3_1674 = address_decode_4(addr_selector2_104[10],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1674,addr_remain3_1674);


wire[15:0] addr_selector3_1675;
wire[15:0] addr_remain3_1675;
address_decode_4 decoder_3_1675 = address_decode_4(addr_selector2_104[11],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1675,addr_remain3_1675);


wire[15:0] addr_selector3_1676;
wire[15:0] addr_remain3_1676;
address_decode_4 decoder_3_1676 = address_decode_4(addr_selector2_104[12],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1676,addr_remain3_1676);


wire[15:0] addr_selector3_1677;
wire[15:0] addr_remain3_1677;
address_decode_4 decoder_3_1677 = address_decode_4(addr_selector2_104[13],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1677,addr_remain3_1677);


wire[15:0] addr_selector3_1678;
wire[15:0] addr_remain3_1678;
address_decode_4 decoder_3_1678 = address_decode_4(addr_selector2_104[14],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1678,addr_remain3_1678);


wire[15:0] addr_selector3_1679;
wire[15:0] addr_remain3_1679;
address_decode_4 decoder_3_1679 = address_decode_4(addr_selector2_104[15],addr_remain2_104[15:0],addr_remain2_104,addr_selector3_1679,addr_remain3_1679);


wire[15:0] addr_selector3_1680;
wire[15:0] addr_remain3_1680;
address_decode_4 decoder_3_1680 = address_decode_4(addr_selector2_105[0],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1680,addr_remain3_1680);


wire[15:0] addr_selector3_1681;
wire[15:0] addr_remain3_1681;
address_decode_4 decoder_3_1681 = address_decode_4(addr_selector2_105[1],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1681,addr_remain3_1681);


wire[15:0] addr_selector3_1682;
wire[15:0] addr_remain3_1682;
address_decode_4 decoder_3_1682 = address_decode_4(addr_selector2_105[2],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1682,addr_remain3_1682);


wire[15:0] addr_selector3_1683;
wire[15:0] addr_remain3_1683;
address_decode_4 decoder_3_1683 = address_decode_4(addr_selector2_105[3],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1683,addr_remain3_1683);


wire[15:0] addr_selector3_1684;
wire[15:0] addr_remain3_1684;
address_decode_4 decoder_3_1684 = address_decode_4(addr_selector2_105[4],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1684,addr_remain3_1684);


wire[15:0] addr_selector3_1685;
wire[15:0] addr_remain3_1685;
address_decode_4 decoder_3_1685 = address_decode_4(addr_selector2_105[5],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1685,addr_remain3_1685);


wire[15:0] addr_selector3_1686;
wire[15:0] addr_remain3_1686;
address_decode_4 decoder_3_1686 = address_decode_4(addr_selector2_105[6],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1686,addr_remain3_1686);


wire[15:0] addr_selector3_1687;
wire[15:0] addr_remain3_1687;
address_decode_4 decoder_3_1687 = address_decode_4(addr_selector2_105[7],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1687,addr_remain3_1687);


wire[15:0] addr_selector3_1688;
wire[15:0] addr_remain3_1688;
address_decode_4 decoder_3_1688 = address_decode_4(addr_selector2_105[8],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1688,addr_remain3_1688);


wire[15:0] addr_selector3_1689;
wire[15:0] addr_remain3_1689;
address_decode_4 decoder_3_1689 = address_decode_4(addr_selector2_105[9],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1689,addr_remain3_1689);


wire[15:0] addr_selector3_1690;
wire[15:0] addr_remain3_1690;
address_decode_4 decoder_3_1690 = address_decode_4(addr_selector2_105[10],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1690,addr_remain3_1690);


wire[15:0] addr_selector3_1691;
wire[15:0] addr_remain3_1691;
address_decode_4 decoder_3_1691 = address_decode_4(addr_selector2_105[11],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1691,addr_remain3_1691);


wire[15:0] addr_selector3_1692;
wire[15:0] addr_remain3_1692;
address_decode_4 decoder_3_1692 = address_decode_4(addr_selector2_105[12],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1692,addr_remain3_1692);


wire[15:0] addr_selector3_1693;
wire[15:0] addr_remain3_1693;
address_decode_4 decoder_3_1693 = address_decode_4(addr_selector2_105[13],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1693,addr_remain3_1693);


wire[15:0] addr_selector3_1694;
wire[15:0] addr_remain3_1694;
address_decode_4 decoder_3_1694 = address_decode_4(addr_selector2_105[14],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1694,addr_remain3_1694);


wire[15:0] addr_selector3_1695;
wire[15:0] addr_remain3_1695;
address_decode_4 decoder_3_1695 = address_decode_4(addr_selector2_105[15],addr_remain2_105[15:0],addr_remain2_105,addr_selector3_1695,addr_remain3_1695);


wire[15:0] addr_selector3_1696;
wire[15:0] addr_remain3_1696;
address_decode_4 decoder_3_1696 = address_decode_4(addr_selector2_106[0],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1696,addr_remain3_1696);


wire[15:0] addr_selector3_1697;
wire[15:0] addr_remain3_1697;
address_decode_4 decoder_3_1697 = address_decode_4(addr_selector2_106[1],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1697,addr_remain3_1697);


wire[15:0] addr_selector3_1698;
wire[15:0] addr_remain3_1698;
address_decode_4 decoder_3_1698 = address_decode_4(addr_selector2_106[2],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1698,addr_remain3_1698);


wire[15:0] addr_selector3_1699;
wire[15:0] addr_remain3_1699;
address_decode_4 decoder_3_1699 = address_decode_4(addr_selector2_106[3],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1699,addr_remain3_1699);


wire[15:0] addr_selector3_1700;
wire[15:0] addr_remain3_1700;
address_decode_4 decoder_3_1700 = address_decode_4(addr_selector2_106[4],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1700,addr_remain3_1700);


wire[15:0] addr_selector3_1701;
wire[15:0] addr_remain3_1701;
address_decode_4 decoder_3_1701 = address_decode_4(addr_selector2_106[5],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1701,addr_remain3_1701);


wire[15:0] addr_selector3_1702;
wire[15:0] addr_remain3_1702;
address_decode_4 decoder_3_1702 = address_decode_4(addr_selector2_106[6],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1702,addr_remain3_1702);


wire[15:0] addr_selector3_1703;
wire[15:0] addr_remain3_1703;
address_decode_4 decoder_3_1703 = address_decode_4(addr_selector2_106[7],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1703,addr_remain3_1703);


wire[15:0] addr_selector3_1704;
wire[15:0] addr_remain3_1704;
address_decode_4 decoder_3_1704 = address_decode_4(addr_selector2_106[8],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1704,addr_remain3_1704);


wire[15:0] addr_selector3_1705;
wire[15:0] addr_remain3_1705;
address_decode_4 decoder_3_1705 = address_decode_4(addr_selector2_106[9],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1705,addr_remain3_1705);


wire[15:0] addr_selector3_1706;
wire[15:0] addr_remain3_1706;
address_decode_4 decoder_3_1706 = address_decode_4(addr_selector2_106[10],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1706,addr_remain3_1706);


wire[15:0] addr_selector3_1707;
wire[15:0] addr_remain3_1707;
address_decode_4 decoder_3_1707 = address_decode_4(addr_selector2_106[11],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1707,addr_remain3_1707);


wire[15:0] addr_selector3_1708;
wire[15:0] addr_remain3_1708;
address_decode_4 decoder_3_1708 = address_decode_4(addr_selector2_106[12],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1708,addr_remain3_1708);


wire[15:0] addr_selector3_1709;
wire[15:0] addr_remain3_1709;
address_decode_4 decoder_3_1709 = address_decode_4(addr_selector2_106[13],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1709,addr_remain3_1709);


wire[15:0] addr_selector3_1710;
wire[15:0] addr_remain3_1710;
address_decode_4 decoder_3_1710 = address_decode_4(addr_selector2_106[14],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1710,addr_remain3_1710);


wire[15:0] addr_selector3_1711;
wire[15:0] addr_remain3_1711;
address_decode_4 decoder_3_1711 = address_decode_4(addr_selector2_106[15],addr_remain2_106[15:0],addr_remain2_106,addr_selector3_1711,addr_remain3_1711);


wire[15:0] addr_selector3_1712;
wire[15:0] addr_remain3_1712;
address_decode_4 decoder_3_1712 = address_decode_4(addr_selector2_107[0],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1712,addr_remain3_1712);


wire[15:0] addr_selector3_1713;
wire[15:0] addr_remain3_1713;
address_decode_4 decoder_3_1713 = address_decode_4(addr_selector2_107[1],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1713,addr_remain3_1713);


wire[15:0] addr_selector3_1714;
wire[15:0] addr_remain3_1714;
address_decode_4 decoder_3_1714 = address_decode_4(addr_selector2_107[2],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1714,addr_remain3_1714);


wire[15:0] addr_selector3_1715;
wire[15:0] addr_remain3_1715;
address_decode_4 decoder_3_1715 = address_decode_4(addr_selector2_107[3],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1715,addr_remain3_1715);


wire[15:0] addr_selector3_1716;
wire[15:0] addr_remain3_1716;
address_decode_4 decoder_3_1716 = address_decode_4(addr_selector2_107[4],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1716,addr_remain3_1716);


wire[15:0] addr_selector3_1717;
wire[15:0] addr_remain3_1717;
address_decode_4 decoder_3_1717 = address_decode_4(addr_selector2_107[5],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1717,addr_remain3_1717);


wire[15:0] addr_selector3_1718;
wire[15:0] addr_remain3_1718;
address_decode_4 decoder_3_1718 = address_decode_4(addr_selector2_107[6],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1718,addr_remain3_1718);


wire[15:0] addr_selector3_1719;
wire[15:0] addr_remain3_1719;
address_decode_4 decoder_3_1719 = address_decode_4(addr_selector2_107[7],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1719,addr_remain3_1719);


wire[15:0] addr_selector3_1720;
wire[15:0] addr_remain3_1720;
address_decode_4 decoder_3_1720 = address_decode_4(addr_selector2_107[8],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1720,addr_remain3_1720);


wire[15:0] addr_selector3_1721;
wire[15:0] addr_remain3_1721;
address_decode_4 decoder_3_1721 = address_decode_4(addr_selector2_107[9],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1721,addr_remain3_1721);


wire[15:0] addr_selector3_1722;
wire[15:0] addr_remain3_1722;
address_decode_4 decoder_3_1722 = address_decode_4(addr_selector2_107[10],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1722,addr_remain3_1722);


wire[15:0] addr_selector3_1723;
wire[15:0] addr_remain3_1723;
address_decode_4 decoder_3_1723 = address_decode_4(addr_selector2_107[11],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1723,addr_remain3_1723);


wire[15:0] addr_selector3_1724;
wire[15:0] addr_remain3_1724;
address_decode_4 decoder_3_1724 = address_decode_4(addr_selector2_107[12],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1724,addr_remain3_1724);


wire[15:0] addr_selector3_1725;
wire[15:0] addr_remain3_1725;
address_decode_4 decoder_3_1725 = address_decode_4(addr_selector2_107[13],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1725,addr_remain3_1725);


wire[15:0] addr_selector3_1726;
wire[15:0] addr_remain3_1726;
address_decode_4 decoder_3_1726 = address_decode_4(addr_selector2_107[14],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1726,addr_remain3_1726);


wire[15:0] addr_selector3_1727;
wire[15:0] addr_remain3_1727;
address_decode_4 decoder_3_1727 = address_decode_4(addr_selector2_107[15],addr_remain2_107[15:0],addr_remain2_107,addr_selector3_1727,addr_remain3_1727);


wire[15:0] addr_selector3_1728;
wire[15:0] addr_remain3_1728;
address_decode_4 decoder_3_1728 = address_decode_4(addr_selector2_108[0],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1728,addr_remain3_1728);


wire[15:0] addr_selector3_1729;
wire[15:0] addr_remain3_1729;
address_decode_4 decoder_3_1729 = address_decode_4(addr_selector2_108[1],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1729,addr_remain3_1729);


wire[15:0] addr_selector3_1730;
wire[15:0] addr_remain3_1730;
address_decode_4 decoder_3_1730 = address_decode_4(addr_selector2_108[2],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1730,addr_remain3_1730);


wire[15:0] addr_selector3_1731;
wire[15:0] addr_remain3_1731;
address_decode_4 decoder_3_1731 = address_decode_4(addr_selector2_108[3],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1731,addr_remain3_1731);


wire[15:0] addr_selector3_1732;
wire[15:0] addr_remain3_1732;
address_decode_4 decoder_3_1732 = address_decode_4(addr_selector2_108[4],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1732,addr_remain3_1732);


wire[15:0] addr_selector3_1733;
wire[15:0] addr_remain3_1733;
address_decode_4 decoder_3_1733 = address_decode_4(addr_selector2_108[5],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1733,addr_remain3_1733);


wire[15:0] addr_selector3_1734;
wire[15:0] addr_remain3_1734;
address_decode_4 decoder_3_1734 = address_decode_4(addr_selector2_108[6],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1734,addr_remain3_1734);


wire[15:0] addr_selector3_1735;
wire[15:0] addr_remain3_1735;
address_decode_4 decoder_3_1735 = address_decode_4(addr_selector2_108[7],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1735,addr_remain3_1735);


wire[15:0] addr_selector3_1736;
wire[15:0] addr_remain3_1736;
address_decode_4 decoder_3_1736 = address_decode_4(addr_selector2_108[8],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1736,addr_remain3_1736);


wire[15:0] addr_selector3_1737;
wire[15:0] addr_remain3_1737;
address_decode_4 decoder_3_1737 = address_decode_4(addr_selector2_108[9],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1737,addr_remain3_1737);


wire[15:0] addr_selector3_1738;
wire[15:0] addr_remain3_1738;
address_decode_4 decoder_3_1738 = address_decode_4(addr_selector2_108[10],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1738,addr_remain3_1738);


wire[15:0] addr_selector3_1739;
wire[15:0] addr_remain3_1739;
address_decode_4 decoder_3_1739 = address_decode_4(addr_selector2_108[11],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1739,addr_remain3_1739);


wire[15:0] addr_selector3_1740;
wire[15:0] addr_remain3_1740;
address_decode_4 decoder_3_1740 = address_decode_4(addr_selector2_108[12],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1740,addr_remain3_1740);


wire[15:0] addr_selector3_1741;
wire[15:0] addr_remain3_1741;
address_decode_4 decoder_3_1741 = address_decode_4(addr_selector2_108[13],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1741,addr_remain3_1741);


wire[15:0] addr_selector3_1742;
wire[15:0] addr_remain3_1742;
address_decode_4 decoder_3_1742 = address_decode_4(addr_selector2_108[14],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1742,addr_remain3_1742);


wire[15:0] addr_selector3_1743;
wire[15:0] addr_remain3_1743;
address_decode_4 decoder_3_1743 = address_decode_4(addr_selector2_108[15],addr_remain2_108[15:0],addr_remain2_108,addr_selector3_1743,addr_remain3_1743);


wire[15:0] addr_selector3_1744;
wire[15:0] addr_remain3_1744;
address_decode_4 decoder_3_1744 = address_decode_4(addr_selector2_109[0],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1744,addr_remain3_1744);


wire[15:0] addr_selector3_1745;
wire[15:0] addr_remain3_1745;
address_decode_4 decoder_3_1745 = address_decode_4(addr_selector2_109[1],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1745,addr_remain3_1745);


wire[15:0] addr_selector3_1746;
wire[15:0] addr_remain3_1746;
address_decode_4 decoder_3_1746 = address_decode_4(addr_selector2_109[2],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1746,addr_remain3_1746);


wire[15:0] addr_selector3_1747;
wire[15:0] addr_remain3_1747;
address_decode_4 decoder_3_1747 = address_decode_4(addr_selector2_109[3],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1747,addr_remain3_1747);


wire[15:0] addr_selector3_1748;
wire[15:0] addr_remain3_1748;
address_decode_4 decoder_3_1748 = address_decode_4(addr_selector2_109[4],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1748,addr_remain3_1748);


wire[15:0] addr_selector3_1749;
wire[15:0] addr_remain3_1749;
address_decode_4 decoder_3_1749 = address_decode_4(addr_selector2_109[5],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1749,addr_remain3_1749);


wire[15:0] addr_selector3_1750;
wire[15:0] addr_remain3_1750;
address_decode_4 decoder_3_1750 = address_decode_4(addr_selector2_109[6],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1750,addr_remain3_1750);


wire[15:0] addr_selector3_1751;
wire[15:0] addr_remain3_1751;
address_decode_4 decoder_3_1751 = address_decode_4(addr_selector2_109[7],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1751,addr_remain3_1751);


wire[15:0] addr_selector3_1752;
wire[15:0] addr_remain3_1752;
address_decode_4 decoder_3_1752 = address_decode_4(addr_selector2_109[8],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1752,addr_remain3_1752);


wire[15:0] addr_selector3_1753;
wire[15:0] addr_remain3_1753;
address_decode_4 decoder_3_1753 = address_decode_4(addr_selector2_109[9],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1753,addr_remain3_1753);


wire[15:0] addr_selector3_1754;
wire[15:0] addr_remain3_1754;
address_decode_4 decoder_3_1754 = address_decode_4(addr_selector2_109[10],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1754,addr_remain3_1754);


wire[15:0] addr_selector3_1755;
wire[15:0] addr_remain3_1755;
address_decode_4 decoder_3_1755 = address_decode_4(addr_selector2_109[11],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1755,addr_remain3_1755);


wire[15:0] addr_selector3_1756;
wire[15:0] addr_remain3_1756;
address_decode_4 decoder_3_1756 = address_decode_4(addr_selector2_109[12],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1756,addr_remain3_1756);


wire[15:0] addr_selector3_1757;
wire[15:0] addr_remain3_1757;
address_decode_4 decoder_3_1757 = address_decode_4(addr_selector2_109[13],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1757,addr_remain3_1757);


wire[15:0] addr_selector3_1758;
wire[15:0] addr_remain3_1758;
address_decode_4 decoder_3_1758 = address_decode_4(addr_selector2_109[14],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1758,addr_remain3_1758);


wire[15:0] addr_selector3_1759;
wire[15:0] addr_remain3_1759;
address_decode_4 decoder_3_1759 = address_decode_4(addr_selector2_109[15],addr_remain2_109[15:0],addr_remain2_109,addr_selector3_1759,addr_remain3_1759);


wire[15:0] addr_selector3_1760;
wire[15:0] addr_remain3_1760;
address_decode_4 decoder_3_1760 = address_decode_4(addr_selector2_110[0],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1760,addr_remain3_1760);


wire[15:0] addr_selector3_1761;
wire[15:0] addr_remain3_1761;
address_decode_4 decoder_3_1761 = address_decode_4(addr_selector2_110[1],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1761,addr_remain3_1761);


wire[15:0] addr_selector3_1762;
wire[15:0] addr_remain3_1762;
address_decode_4 decoder_3_1762 = address_decode_4(addr_selector2_110[2],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1762,addr_remain3_1762);


wire[15:0] addr_selector3_1763;
wire[15:0] addr_remain3_1763;
address_decode_4 decoder_3_1763 = address_decode_4(addr_selector2_110[3],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1763,addr_remain3_1763);


wire[15:0] addr_selector3_1764;
wire[15:0] addr_remain3_1764;
address_decode_4 decoder_3_1764 = address_decode_4(addr_selector2_110[4],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1764,addr_remain3_1764);


wire[15:0] addr_selector3_1765;
wire[15:0] addr_remain3_1765;
address_decode_4 decoder_3_1765 = address_decode_4(addr_selector2_110[5],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1765,addr_remain3_1765);


wire[15:0] addr_selector3_1766;
wire[15:0] addr_remain3_1766;
address_decode_4 decoder_3_1766 = address_decode_4(addr_selector2_110[6],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1766,addr_remain3_1766);


wire[15:0] addr_selector3_1767;
wire[15:0] addr_remain3_1767;
address_decode_4 decoder_3_1767 = address_decode_4(addr_selector2_110[7],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1767,addr_remain3_1767);


wire[15:0] addr_selector3_1768;
wire[15:0] addr_remain3_1768;
address_decode_4 decoder_3_1768 = address_decode_4(addr_selector2_110[8],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1768,addr_remain3_1768);


wire[15:0] addr_selector3_1769;
wire[15:0] addr_remain3_1769;
address_decode_4 decoder_3_1769 = address_decode_4(addr_selector2_110[9],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1769,addr_remain3_1769);


wire[15:0] addr_selector3_1770;
wire[15:0] addr_remain3_1770;
address_decode_4 decoder_3_1770 = address_decode_4(addr_selector2_110[10],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1770,addr_remain3_1770);


wire[15:0] addr_selector3_1771;
wire[15:0] addr_remain3_1771;
address_decode_4 decoder_3_1771 = address_decode_4(addr_selector2_110[11],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1771,addr_remain3_1771);


wire[15:0] addr_selector3_1772;
wire[15:0] addr_remain3_1772;
address_decode_4 decoder_3_1772 = address_decode_4(addr_selector2_110[12],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1772,addr_remain3_1772);


wire[15:0] addr_selector3_1773;
wire[15:0] addr_remain3_1773;
address_decode_4 decoder_3_1773 = address_decode_4(addr_selector2_110[13],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1773,addr_remain3_1773);


wire[15:0] addr_selector3_1774;
wire[15:0] addr_remain3_1774;
address_decode_4 decoder_3_1774 = address_decode_4(addr_selector2_110[14],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1774,addr_remain3_1774);


wire[15:0] addr_selector3_1775;
wire[15:0] addr_remain3_1775;
address_decode_4 decoder_3_1775 = address_decode_4(addr_selector2_110[15],addr_remain2_110[15:0],addr_remain2_110,addr_selector3_1775,addr_remain3_1775);


wire[15:0] addr_selector3_1776;
wire[15:0] addr_remain3_1776;
address_decode_4 decoder_3_1776 = address_decode_4(addr_selector2_111[0],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1776,addr_remain3_1776);


wire[15:0] addr_selector3_1777;
wire[15:0] addr_remain3_1777;
address_decode_4 decoder_3_1777 = address_decode_4(addr_selector2_111[1],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1777,addr_remain3_1777);


wire[15:0] addr_selector3_1778;
wire[15:0] addr_remain3_1778;
address_decode_4 decoder_3_1778 = address_decode_4(addr_selector2_111[2],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1778,addr_remain3_1778);


wire[15:0] addr_selector3_1779;
wire[15:0] addr_remain3_1779;
address_decode_4 decoder_3_1779 = address_decode_4(addr_selector2_111[3],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1779,addr_remain3_1779);


wire[15:0] addr_selector3_1780;
wire[15:0] addr_remain3_1780;
address_decode_4 decoder_3_1780 = address_decode_4(addr_selector2_111[4],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1780,addr_remain3_1780);


wire[15:0] addr_selector3_1781;
wire[15:0] addr_remain3_1781;
address_decode_4 decoder_3_1781 = address_decode_4(addr_selector2_111[5],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1781,addr_remain3_1781);


wire[15:0] addr_selector3_1782;
wire[15:0] addr_remain3_1782;
address_decode_4 decoder_3_1782 = address_decode_4(addr_selector2_111[6],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1782,addr_remain3_1782);


wire[15:0] addr_selector3_1783;
wire[15:0] addr_remain3_1783;
address_decode_4 decoder_3_1783 = address_decode_4(addr_selector2_111[7],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1783,addr_remain3_1783);


wire[15:0] addr_selector3_1784;
wire[15:0] addr_remain3_1784;
address_decode_4 decoder_3_1784 = address_decode_4(addr_selector2_111[8],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1784,addr_remain3_1784);


wire[15:0] addr_selector3_1785;
wire[15:0] addr_remain3_1785;
address_decode_4 decoder_3_1785 = address_decode_4(addr_selector2_111[9],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1785,addr_remain3_1785);


wire[15:0] addr_selector3_1786;
wire[15:0] addr_remain3_1786;
address_decode_4 decoder_3_1786 = address_decode_4(addr_selector2_111[10],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1786,addr_remain3_1786);


wire[15:0] addr_selector3_1787;
wire[15:0] addr_remain3_1787;
address_decode_4 decoder_3_1787 = address_decode_4(addr_selector2_111[11],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1787,addr_remain3_1787);


wire[15:0] addr_selector3_1788;
wire[15:0] addr_remain3_1788;
address_decode_4 decoder_3_1788 = address_decode_4(addr_selector2_111[12],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1788,addr_remain3_1788);


wire[15:0] addr_selector3_1789;
wire[15:0] addr_remain3_1789;
address_decode_4 decoder_3_1789 = address_decode_4(addr_selector2_111[13],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1789,addr_remain3_1789);


wire[15:0] addr_selector3_1790;
wire[15:0] addr_remain3_1790;
address_decode_4 decoder_3_1790 = address_decode_4(addr_selector2_111[14],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1790,addr_remain3_1790);


wire[15:0] addr_selector3_1791;
wire[15:0] addr_remain3_1791;
address_decode_4 decoder_3_1791 = address_decode_4(addr_selector2_111[15],addr_remain2_111[15:0],addr_remain2_111,addr_selector3_1791,addr_remain3_1791);


wire[15:0] addr_selector3_1792;
wire[15:0] addr_remain3_1792;
address_decode_4 decoder_3_1792 = address_decode_4(addr_selector2_112[0],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1792,addr_remain3_1792);


wire[15:0] addr_selector3_1793;
wire[15:0] addr_remain3_1793;
address_decode_4 decoder_3_1793 = address_decode_4(addr_selector2_112[1],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1793,addr_remain3_1793);


wire[15:0] addr_selector3_1794;
wire[15:0] addr_remain3_1794;
address_decode_4 decoder_3_1794 = address_decode_4(addr_selector2_112[2],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1794,addr_remain3_1794);


wire[15:0] addr_selector3_1795;
wire[15:0] addr_remain3_1795;
address_decode_4 decoder_3_1795 = address_decode_4(addr_selector2_112[3],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1795,addr_remain3_1795);


wire[15:0] addr_selector3_1796;
wire[15:0] addr_remain3_1796;
address_decode_4 decoder_3_1796 = address_decode_4(addr_selector2_112[4],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1796,addr_remain3_1796);


wire[15:0] addr_selector3_1797;
wire[15:0] addr_remain3_1797;
address_decode_4 decoder_3_1797 = address_decode_4(addr_selector2_112[5],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1797,addr_remain3_1797);


wire[15:0] addr_selector3_1798;
wire[15:0] addr_remain3_1798;
address_decode_4 decoder_3_1798 = address_decode_4(addr_selector2_112[6],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1798,addr_remain3_1798);


wire[15:0] addr_selector3_1799;
wire[15:0] addr_remain3_1799;
address_decode_4 decoder_3_1799 = address_decode_4(addr_selector2_112[7],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1799,addr_remain3_1799);


wire[15:0] addr_selector3_1800;
wire[15:0] addr_remain3_1800;
address_decode_4 decoder_3_1800 = address_decode_4(addr_selector2_112[8],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1800,addr_remain3_1800);


wire[15:0] addr_selector3_1801;
wire[15:0] addr_remain3_1801;
address_decode_4 decoder_3_1801 = address_decode_4(addr_selector2_112[9],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1801,addr_remain3_1801);


wire[15:0] addr_selector3_1802;
wire[15:0] addr_remain3_1802;
address_decode_4 decoder_3_1802 = address_decode_4(addr_selector2_112[10],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1802,addr_remain3_1802);


wire[15:0] addr_selector3_1803;
wire[15:0] addr_remain3_1803;
address_decode_4 decoder_3_1803 = address_decode_4(addr_selector2_112[11],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1803,addr_remain3_1803);


wire[15:0] addr_selector3_1804;
wire[15:0] addr_remain3_1804;
address_decode_4 decoder_3_1804 = address_decode_4(addr_selector2_112[12],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1804,addr_remain3_1804);


wire[15:0] addr_selector3_1805;
wire[15:0] addr_remain3_1805;
address_decode_4 decoder_3_1805 = address_decode_4(addr_selector2_112[13],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1805,addr_remain3_1805);


wire[15:0] addr_selector3_1806;
wire[15:0] addr_remain3_1806;
address_decode_4 decoder_3_1806 = address_decode_4(addr_selector2_112[14],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1806,addr_remain3_1806);


wire[15:0] addr_selector3_1807;
wire[15:0] addr_remain3_1807;
address_decode_4 decoder_3_1807 = address_decode_4(addr_selector2_112[15],addr_remain2_112[15:0],addr_remain2_112,addr_selector3_1807,addr_remain3_1807);


wire[15:0] addr_selector3_1808;
wire[15:0] addr_remain3_1808;
address_decode_4 decoder_3_1808 = address_decode_4(addr_selector2_113[0],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1808,addr_remain3_1808);


wire[15:0] addr_selector3_1809;
wire[15:0] addr_remain3_1809;
address_decode_4 decoder_3_1809 = address_decode_4(addr_selector2_113[1],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1809,addr_remain3_1809);


wire[15:0] addr_selector3_1810;
wire[15:0] addr_remain3_1810;
address_decode_4 decoder_3_1810 = address_decode_4(addr_selector2_113[2],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1810,addr_remain3_1810);


wire[15:0] addr_selector3_1811;
wire[15:0] addr_remain3_1811;
address_decode_4 decoder_3_1811 = address_decode_4(addr_selector2_113[3],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1811,addr_remain3_1811);


wire[15:0] addr_selector3_1812;
wire[15:0] addr_remain3_1812;
address_decode_4 decoder_3_1812 = address_decode_4(addr_selector2_113[4],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1812,addr_remain3_1812);


wire[15:0] addr_selector3_1813;
wire[15:0] addr_remain3_1813;
address_decode_4 decoder_3_1813 = address_decode_4(addr_selector2_113[5],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1813,addr_remain3_1813);


wire[15:0] addr_selector3_1814;
wire[15:0] addr_remain3_1814;
address_decode_4 decoder_3_1814 = address_decode_4(addr_selector2_113[6],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1814,addr_remain3_1814);


wire[15:0] addr_selector3_1815;
wire[15:0] addr_remain3_1815;
address_decode_4 decoder_3_1815 = address_decode_4(addr_selector2_113[7],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1815,addr_remain3_1815);


wire[15:0] addr_selector3_1816;
wire[15:0] addr_remain3_1816;
address_decode_4 decoder_3_1816 = address_decode_4(addr_selector2_113[8],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1816,addr_remain3_1816);


wire[15:0] addr_selector3_1817;
wire[15:0] addr_remain3_1817;
address_decode_4 decoder_3_1817 = address_decode_4(addr_selector2_113[9],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1817,addr_remain3_1817);


wire[15:0] addr_selector3_1818;
wire[15:0] addr_remain3_1818;
address_decode_4 decoder_3_1818 = address_decode_4(addr_selector2_113[10],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1818,addr_remain3_1818);


wire[15:0] addr_selector3_1819;
wire[15:0] addr_remain3_1819;
address_decode_4 decoder_3_1819 = address_decode_4(addr_selector2_113[11],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1819,addr_remain3_1819);


wire[15:0] addr_selector3_1820;
wire[15:0] addr_remain3_1820;
address_decode_4 decoder_3_1820 = address_decode_4(addr_selector2_113[12],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1820,addr_remain3_1820);


wire[15:0] addr_selector3_1821;
wire[15:0] addr_remain3_1821;
address_decode_4 decoder_3_1821 = address_decode_4(addr_selector2_113[13],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1821,addr_remain3_1821);


wire[15:0] addr_selector3_1822;
wire[15:0] addr_remain3_1822;
address_decode_4 decoder_3_1822 = address_decode_4(addr_selector2_113[14],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1822,addr_remain3_1822);


wire[15:0] addr_selector3_1823;
wire[15:0] addr_remain3_1823;
address_decode_4 decoder_3_1823 = address_decode_4(addr_selector2_113[15],addr_remain2_113[15:0],addr_remain2_113,addr_selector3_1823,addr_remain3_1823);


wire[15:0] addr_selector3_1824;
wire[15:0] addr_remain3_1824;
address_decode_4 decoder_3_1824 = address_decode_4(addr_selector2_114[0],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1824,addr_remain3_1824);


wire[15:0] addr_selector3_1825;
wire[15:0] addr_remain3_1825;
address_decode_4 decoder_3_1825 = address_decode_4(addr_selector2_114[1],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1825,addr_remain3_1825);


wire[15:0] addr_selector3_1826;
wire[15:0] addr_remain3_1826;
address_decode_4 decoder_3_1826 = address_decode_4(addr_selector2_114[2],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1826,addr_remain3_1826);


wire[15:0] addr_selector3_1827;
wire[15:0] addr_remain3_1827;
address_decode_4 decoder_3_1827 = address_decode_4(addr_selector2_114[3],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1827,addr_remain3_1827);


wire[15:0] addr_selector3_1828;
wire[15:0] addr_remain3_1828;
address_decode_4 decoder_3_1828 = address_decode_4(addr_selector2_114[4],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1828,addr_remain3_1828);


wire[15:0] addr_selector3_1829;
wire[15:0] addr_remain3_1829;
address_decode_4 decoder_3_1829 = address_decode_4(addr_selector2_114[5],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1829,addr_remain3_1829);


wire[15:0] addr_selector3_1830;
wire[15:0] addr_remain3_1830;
address_decode_4 decoder_3_1830 = address_decode_4(addr_selector2_114[6],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1830,addr_remain3_1830);


wire[15:0] addr_selector3_1831;
wire[15:0] addr_remain3_1831;
address_decode_4 decoder_3_1831 = address_decode_4(addr_selector2_114[7],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1831,addr_remain3_1831);


wire[15:0] addr_selector3_1832;
wire[15:0] addr_remain3_1832;
address_decode_4 decoder_3_1832 = address_decode_4(addr_selector2_114[8],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1832,addr_remain3_1832);


wire[15:0] addr_selector3_1833;
wire[15:0] addr_remain3_1833;
address_decode_4 decoder_3_1833 = address_decode_4(addr_selector2_114[9],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1833,addr_remain3_1833);


wire[15:0] addr_selector3_1834;
wire[15:0] addr_remain3_1834;
address_decode_4 decoder_3_1834 = address_decode_4(addr_selector2_114[10],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1834,addr_remain3_1834);


wire[15:0] addr_selector3_1835;
wire[15:0] addr_remain3_1835;
address_decode_4 decoder_3_1835 = address_decode_4(addr_selector2_114[11],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1835,addr_remain3_1835);


wire[15:0] addr_selector3_1836;
wire[15:0] addr_remain3_1836;
address_decode_4 decoder_3_1836 = address_decode_4(addr_selector2_114[12],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1836,addr_remain3_1836);


wire[15:0] addr_selector3_1837;
wire[15:0] addr_remain3_1837;
address_decode_4 decoder_3_1837 = address_decode_4(addr_selector2_114[13],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1837,addr_remain3_1837);


wire[15:0] addr_selector3_1838;
wire[15:0] addr_remain3_1838;
address_decode_4 decoder_3_1838 = address_decode_4(addr_selector2_114[14],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1838,addr_remain3_1838);


wire[15:0] addr_selector3_1839;
wire[15:0] addr_remain3_1839;
address_decode_4 decoder_3_1839 = address_decode_4(addr_selector2_114[15],addr_remain2_114[15:0],addr_remain2_114,addr_selector3_1839,addr_remain3_1839);


wire[15:0] addr_selector3_1840;
wire[15:0] addr_remain3_1840;
address_decode_4 decoder_3_1840 = address_decode_4(addr_selector2_115[0],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1840,addr_remain3_1840);


wire[15:0] addr_selector3_1841;
wire[15:0] addr_remain3_1841;
address_decode_4 decoder_3_1841 = address_decode_4(addr_selector2_115[1],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1841,addr_remain3_1841);


wire[15:0] addr_selector3_1842;
wire[15:0] addr_remain3_1842;
address_decode_4 decoder_3_1842 = address_decode_4(addr_selector2_115[2],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1842,addr_remain3_1842);


wire[15:0] addr_selector3_1843;
wire[15:0] addr_remain3_1843;
address_decode_4 decoder_3_1843 = address_decode_4(addr_selector2_115[3],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1843,addr_remain3_1843);


wire[15:0] addr_selector3_1844;
wire[15:0] addr_remain3_1844;
address_decode_4 decoder_3_1844 = address_decode_4(addr_selector2_115[4],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1844,addr_remain3_1844);


wire[15:0] addr_selector3_1845;
wire[15:0] addr_remain3_1845;
address_decode_4 decoder_3_1845 = address_decode_4(addr_selector2_115[5],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1845,addr_remain3_1845);


wire[15:0] addr_selector3_1846;
wire[15:0] addr_remain3_1846;
address_decode_4 decoder_3_1846 = address_decode_4(addr_selector2_115[6],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1846,addr_remain3_1846);


wire[15:0] addr_selector3_1847;
wire[15:0] addr_remain3_1847;
address_decode_4 decoder_3_1847 = address_decode_4(addr_selector2_115[7],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1847,addr_remain3_1847);


wire[15:0] addr_selector3_1848;
wire[15:0] addr_remain3_1848;
address_decode_4 decoder_3_1848 = address_decode_4(addr_selector2_115[8],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1848,addr_remain3_1848);


wire[15:0] addr_selector3_1849;
wire[15:0] addr_remain3_1849;
address_decode_4 decoder_3_1849 = address_decode_4(addr_selector2_115[9],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1849,addr_remain3_1849);


wire[15:0] addr_selector3_1850;
wire[15:0] addr_remain3_1850;
address_decode_4 decoder_3_1850 = address_decode_4(addr_selector2_115[10],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1850,addr_remain3_1850);


wire[15:0] addr_selector3_1851;
wire[15:0] addr_remain3_1851;
address_decode_4 decoder_3_1851 = address_decode_4(addr_selector2_115[11],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1851,addr_remain3_1851);


wire[15:0] addr_selector3_1852;
wire[15:0] addr_remain3_1852;
address_decode_4 decoder_3_1852 = address_decode_4(addr_selector2_115[12],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1852,addr_remain3_1852);


wire[15:0] addr_selector3_1853;
wire[15:0] addr_remain3_1853;
address_decode_4 decoder_3_1853 = address_decode_4(addr_selector2_115[13],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1853,addr_remain3_1853);


wire[15:0] addr_selector3_1854;
wire[15:0] addr_remain3_1854;
address_decode_4 decoder_3_1854 = address_decode_4(addr_selector2_115[14],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1854,addr_remain3_1854);


wire[15:0] addr_selector3_1855;
wire[15:0] addr_remain3_1855;
address_decode_4 decoder_3_1855 = address_decode_4(addr_selector2_115[15],addr_remain2_115[15:0],addr_remain2_115,addr_selector3_1855,addr_remain3_1855);


wire[15:0] addr_selector3_1856;
wire[15:0] addr_remain3_1856;
address_decode_4 decoder_3_1856 = address_decode_4(addr_selector2_116[0],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1856,addr_remain3_1856);


wire[15:0] addr_selector3_1857;
wire[15:0] addr_remain3_1857;
address_decode_4 decoder_3_1857 = address_decode_4(addr_selector2_116[1],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1857,addr_remain3_1857);


wire[15:0] addr_selector3_1858;
wire[15:0] addr_remain3_1858;
address_decode_4 decoder_3_1858 = address_decode_4(addr_selector2_116[2],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1858,addr_remain3_1858);


wire[15:0] addr_selector3_1859;
wire[15:0] addr_remain3_1859;
address_decode_4 decoder_3_1859 = address_decode_4(addr_selector2_116[3],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1859,addr_remain3_1859);


wire[15:0] addr_selector3_1860;
wire[15:0] addr_remain3_1860;
address_decode_4 decoder_3_1860 = address_decode_4(addr_selector2_116[4],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1860,addr_remain3_1860);


wire[15:0] addr_selector3_1861;
wire[15:0] addr_remain3_1861;
address_decode_4 decoder_3_1861 = address_decode_4(addr_selector2_116[5],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1861,addr_remain3_1861);


wire[15:0] addr_selector3_1862;
wire[15:0] addr_remain3_1862;
address_decode_4 decoder_3_1862 = address_decode_4(addr_selector2_116[6],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1862,addr_remain3_1862);


wire[15:0] addr_selector3_1863;
wire[15:0] addr_remain3_1863;
address_decode_4 decoder_3_1863 = address_decode_4(addr_selector2_116[7],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1863,addr_remain3_1863);


wire[15:0] addr_selector3_1864;
wire[15:0] addr_remain3_1864;
address_decode_4 decoder_3_1864 = address_decode_4(addr_selector2_116[8],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1864,addr_remain3_1864);


wire[15:0] addr_selector3_1865;
wire[15:0] addr_remain3_1865;
address_decode_4 decoder_3_1865 = address_decode_4(addr_selector2_116[9],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1865,addr_remain3_1865);


wire[15:0] addr_selector3_1866;
wire[15:0] addr_remain3_1866;
address_decode_4 decoder_3_1866 = address_decode_4(addr_selector2_116[10],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1866,addr_remain3_1866);


wire[15:0] addr_selector3_1867;
wire[15:0] addr_remain3_1867;
address_decode_4 decoder_3_1867 = address_decode_4(addr_selector2_116[11],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1867,addr_remain3_1867);


wire[15:0] addr_selector3_1868;
wire[15:0] addr_remain3_1868;
address_decode_4 decoder_3_1868 = address_decode_4(addr_selector2_116[12],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1868,addr_remain3_1868);


wire[15:0] addr_selector3_1869;
wire[15:0] addr_remain3_1869;
address_decode_4 decoder_3_1869 = address_decode_4(addr_selector2_116[13],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1869,addr_remain3_1869);


wire[15:0] addr_selector3_1870;
wire[15:0] addr_remain3_1870;
address_decode_4 decoder_3_1870 = address_decode_4(addr_selector2_116[14],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1870,addr_remain3_1870);


wire[15:0] addr_selector3_1871;
wire[15:0] addr_remain3_1871;
address_decode_4 decoder_3_1871 = address_decode_4(addr_selector2_116[15],addr_remain2_116[15:0],addr_remain2_116,addr_selector3_1871,addr_remain3_1871);


wire[15:0] addr_selector3_1872;
wire[15:0] addr_remain3_1872;
address_decode_4 decoder_3_1872 = address_decode_4(addr_selector2_117[0],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1872,addr_remain3_1872);


wire[15:0] addr_selector3_1873;
wire[15:0] addr_remain3_1873;
address_decode_4 decoder_3_1873 = address_decode_4(addr_selector2_117[1],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1873,addr_remain3_1873);


wire[15:0] addr_selector3_1874;
wire[15:0] addr_remain3_1874;
address_decode_4 decoder_3_1874 = address_decode_4(addr_selector2_117[2],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1874,addr_remain3_1874);


wire[15:0] addr_selector3_1875;
wire[15:0] addr_remain3_1875;
address_decode_4 decoder_3_1875 = address_decode_4(addr_selector2_117[3],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1875,addr_remain3_1875);


wire[15:0] addr_selector3_1876;
wire[15:0] addr_remain3_1876;
address_decode_4 decoder_3_1876 = address_decode_4(addr_selector2_117[4],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1876,addr_remain3_1876);


wire[15:0] addr_selector3_1877;
wire[15:0] addr_remain3_1877;
address_decode_4 decoder_3_1877 = address_decode_4(addr_selector2_117[5],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1877,addr_remain3_1877);


wire[15:0] addr_selector3_1878;
wire[15:0] addr_remain3_1878;
address_decode_4 decoder_3_1878 = address_decode_4(addr_selector2_117[6],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1878,addr_remain3_1878);


wire[15:0] addr_selector3_1879;
wire[15:0] addr_remain3_1879;
address_decode_4 decoder_3_1879 = address_decode_4(addr_selector2_117[7],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1879,addr_remain3_1879);


wire[15:0] addr_selector3_1880;
wire[15:0] addr_remain3_1880;
address_decode_4 decoder_3_1880 = address_decode_4(addr_selector2_117[8],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1880,addr_remain3_1880);


wire[15:0] addr_selector3_1881;
wire[15:0] addr_remain3_1881;
address_decode_4 decoder_3_1881 = address_decode_4(addr_selector2_117[9],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1881,addr_remain3_1881);


wire[15:0] addr_selector3_1882;
wire[15:0] addr_remain3_1882;
address_decode_4 decoder_3_1882 = address_decode_4(addr_selector2_117[10],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1882,addr_remain3_1882);


wire[15:0] addr_selector3_1883;
wire[15:0] addr_remain3_1883;
address_decode_4 decoder_3_1883 = address_decode_4(addr_selector2_117[11],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1883,addr_remain3_1883);


wire[15:0] addr_selector3_1884;
wire[15:0] addr_remain3_1884;
address_decode_4 decoder_3_1884 = address_decode_4(addr_selector2_117[12],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1884,addr_remain3_1884);


wire[15:0] addr_selector3_1885;
wire[15:0] addr_remain3_1885;
address_decode_4 decoder_3_1885 = address_decode_4(addr_selector2_117[13],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1885,addr_remain3_1885);


wire[15:0] addr_selector3_1886;
wire[15:0] addr_remain3_1886;
address_decode_4 decoder_3_1886 = address_decode_4(addr_selector2_117[14],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1886,addr_remain3_1886);


wire[15:0] addr_selector3_1887;
wire[15:0] addr_remain3_1887;
address_decode_4 decoder_3_1887 = address_decode_4(addr_selector2_117[15],addr_remain2_117[15:0],addr_remain2_117,addr_selector3_1887,addr_remain3_1887);


wire[15:0] addr_selector3_1888;
wire[15:0] addr_remain3_1888;
address_decode_4 decoder_3_1888 = address_decode_4(addr_selector2_118[0],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1888,addr_remain3_1888);


wire[15:0] addr_selector3_1889;
wire[15:0] addr_remain3_1889;
address_decode_4 decoder_3_1889 = address_decode_4(addr_selector2_118[1],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1889,addr_remain3_1889);


wire[15:0] addr_selector3_1890;
wire[15:0] addr_remain3_1890;
address_decode_4 decoder_3_1890 = address_decode_4(addr_selector2_118[2],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1890,addr_remain3_1890);


wire[15:0] addr_selector3_1891;
wire[15:0] addr_remain3_1891;
address_decode_4 decoder_3_1891 = address_decode_4(addr_selector2_118[3],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1891,addr_remain3_1891);


wire[15:0] addr_selector3_1892;
wire[15:0] addr_remain3_1892;
address_decode_4 decoder_3_1892 = address_decode_4(addr_selector2_118[4],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1892,addr_remain3_1892);


wire[15:0] addr_selector3_1893;
wire[15:0] addr_remain3_1893;
address_decode_4 decoder_3_1893 = address_decode_4(addr_selector2_118[5],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1893,addr_remain3_1893);


wire[15:0] addr_selector3_1894;
wire[15:0] addr_remain3_1894;
address_decode_4 decoder_3_1894 = address_decode_4(addr_selector2_118[6],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1894,addr_remain3_1894);


wire[15:0] addr_selector3_1895;
wire[15:0] addr_remain3_1895;
address_decode_4 decoder_3_1895 = address_decode_4(addr_selector2_118[7],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1895,addr_remain3_1895);


wire[15:0] addr_selector3_1896;
wire[15:0] addr_remain3_1896;
address_decode_4 decoder_3_1896 = address_decode_4(addr_selector2_118[8],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1896,addr_remain3_1896);


wire[15:0] addr_selector3_1897;
wire[15:0] addr_remain3_1897;
address_decode_4 decoder_3_1897 = address_decode_4(addr_selector2_118[9],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1897,addr_remain3_1897);


wire[15:0] addr_selector3_1898;
wire[15:0] addr_remain3_1898;
address_decode_4 decoder_3_1898 = address_decode_4(addr_selector2_118[10],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1898,addr_remain3_1898);


wire[15:0] addr_selector3_1899;
wire[15:0] addr_remain3_1899;
address_decode_4 decoder_3_1899 = address_decode_4(addr_selector2_118[11],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1899,addr_remain3_1899);


wire[15:0] addr_selector3_1900;
wire[15:0] addr_remain3_1900;
address_decode_4 decoder_3_1900 = address_decode_4(addr_selector2_118[12],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1900,addr_remain3_1900);


wire[15:0] addr_selector3_1901;
wire[15:0] addr_remain3_1901;
address_decode_4 decoder_3_1901 = address_decode_4(addr_selector2_118[13],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1901,addr_remain3_1901);


wire[15:0] addr_selector3_1902;
wire[15:0] addr_remain3_1902;
address_decode_4 decoder_3_1902 = address_decode_4(addr_selector2_118[14],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1902,addr_remain3_1902);


wire[15:0] addr_selector3_1903;
wire[15:0] addr_remain3_1903;
address_decode_4 decoder_3_1903 = address_decode_4(addr_selector2_118[15],addr_remain2_118[15:0],addr_remain2_118,addr_selector3_1903,addr_remain3_1903);


wire[15:0] addr_selector3_1904;
wire[15:0] addr_remain3_1904;
address_decode_4 decoder_3_1904 = address_decode_4(addr_selector2_119[0],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1904,addr_remain3_1904);


wire[15:0] addr_selector3_1905;
wire[15:0] addr_remain3_1905;
address_decode_4 decoder_3_1905 = address_decode_4(addr_selector2_119[1],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1905,addr_remain3_1905);


wire[15:0] addr_selector3_1906;
wire[15:0] addr_remain3_1906;
address_decode_4 decoder_3_1906 = address_decode_4(addr_selector2_119[2],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1906,addr_remain3_1906);


wire[15:0] addr_selector3_1907;
wire[15:0] addr_remain3_1907;
address_decode_4 decoder_3_1907 = address_decode_4(addr_selector2_119[3],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1907,addr_remain3_1907);


wire[15:0] addr_selector3_1908;
wire[15:0] addr_remain3_1908;
address_decode_4 decoder_3_1908 = address_decode_4(addr_selector2_119[4],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1908,addr_remain3_1908);


wire[15:0] addr_selector3_1909;
wire[15:0] addr_remain3_1909;
address_decode_4 decoder_3_1909 = address_decode_4(addr_selector2_119[5],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1909,addr_remain3_1909);


wire[15:0] addr_selector3_1910;
wire[15:0] addr_remain3_1910;
address_decode_4 decoder_3_1910 = address_decode_4(addr_selector2_119[6],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1910,addr_remain3_1910);


wire[15:0] addr_selector3_1911;
wire[15:0] addr_remain3_1911;
address_decode_4 decoder_3_1911 = address_decode_4(addr_selector2_119[7],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1911,addr_remain3_1911);


wire[15:0] addr_selector3_1912;
wire[15:0] addr_remain3_1912;
address_decode_4 decoder_3_1912 = address_decode_4(addr_selector2_119[8],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1912,addr_remain3_1912);


wire[15:0] addr_selector3_1913;
wire[15:0] addr_remain3_1913;
address_decode_4 decoder_3_1913 = address_decode_4(addr_selector2_119[9],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1913,addr_remain3_1913);


wire[15:0] addr_selector3_1914;
wire[15:0] addr_remain3_1914;
address_decode_4 decoder_3_1914 = address_decode_4(addr_selector2_119[10],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1914,addr_remain3_1914);


wire[15:0] addr_selector3_1915;
wire[15:0] addr_remain3_1915;
address_decode_4 decoder_3_1915 = address_decode_4(addr_selector2_119[11],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1915,addr_remain3_1915);


wire[15:0] addr_selector3_1916;
wire[15:0] addr_remain3_1916;
address_decode_4 decoder_3_1916 = address_decode_4(addr_selector2_119[12],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1916,addr_remain3_1916);


wire[15:0] addr_selector3_1917;
wire[15:0] addr_remain3_1917;
address_decode_4 decoder_3_1917 = address_decode_4(addr_selector2_119[13],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1917,addr_remain3_1917);


wire[15:0] addr_selector3_1918;
wire[15:0] addr_remain3_1918;
address_decode_4 decoder_3_1918 = address_decode_4(addr_selector2_119[14],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1918,addr_remain3_1918);


wire[15:0] addr_selector3_1919;
wire[15:0] addr_remain3_1919;
address_decode_4 decoder_3_1919 = address_decode_4(addr_selector2_119[15],addr_remain2_119[15:0],addr_remain2_119,addr_selector3_1919,addr_remain3_1919);


wire[15:0] addr_selector3_1920;
wire[15:0] addr_remain3_1920;
address_decode_4 decoder_3_1920 = address_decode_4(addr_selector2_120[0],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1920,addr_remain3_1920);


wire[15:0] addr_selector3_1921;
wire[15:0] addr_remain3_1921;
address_decode_4 decoder_3_1921 = address_decode_4(addr_selector2_120[1],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1921,addr_remain3_1921);


wire[15:0] addr_selector3_1922;
wire[15:0] addr_remain3_1922;
address_decode_4 decoder_3_1922 = address_decode_4(addr_selector2_120[2],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1922,addr_remain3_1922);


wire[15:0] addr_selector3_1923;
wire[15:0] addr_remain3_1923;
address_decode_4 decoder_3_1923 = address_decode_4(addr_selector2_120[3],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1923,addr_remain3_1923);


wire[15:0] addr_selector3_1924;
wire[15:0] addr_remain3_1924;
address_decode_4 decoder_3_1924 = address_decode_4(addr_selector2_120[4],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1924,addr_remain3_1924);


wire[15:0] addr_selector3_1925;
wire[15:0] addr_remain3_1925;
address_decode_4 decoder_3_1925 = address_decode_4(addr_selector2_120[5],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1925,addr_remain3_1925);


wire[15:0] addr_selector3_1926;
wire[15:0] addr_remain3_1926;
address_decode_4 decoder_3_1926 = address_decode_4(addr_selector2_120[6],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1926,addr_remain3_1926);


wire[15:0] addr_selector3_1927;
wire[15:0] addr_remain3_1927;
address_decode_4 decoder_3_1927 = address_decode_4(addr_selector2_120[7],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1927,addr_remain3_1927);


wire[15:0] addr_selector3_1928;
wire[15:0] addr_remain3_1928;
address_decode_4 decoder_3_1928 = address_decode_4(addr_selector2_120[8],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1928,addr_remain3_1928);


wire[15:0] addr_selector3_1929;
wire[15:0] addr_remain3_1929;
address_decode_4 decoder_3_1929 = address_decode_4(addr_selector2_120[9],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1929,addr_remain3_1929);


wire[15:0] addr_selector3_1930;
wire[15:0] addr_remain3_1930;
address_decode_4 decoder_3_1930 = address_decode_4(addr_selector2_120[10],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1930,addr_remain3_1930);


wire[15:0] addr_selector3_1931;
wire[15:0] addr_remain3_1931;
address_decode_4 decoder_3_1931 = address_decode_4(addr_selector2_120[11],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1931,addr_remain3_1931);


wire[15:0] addr_selector3_1932;
wire[15:0] addr_remain3_1932;
address_decode_4 decoder_3_1932 = address_decode_4(addr_selector2_120[12],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1932,addr_remain3_1932);


wire[15:0] addr_selector3_1933;
wire[15:0] addr_remain3_1933;
address_decode_4 decoder_3_1933 = address_decode_4(addr_selector2_120[13],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1933,addr_remain3_1933);


wire[15:0] addr_selector3_1934;
wire[15:0] addr_remain3_1934;
address_decode_4 decoder_3_1934 = address_decode_4(addr_selector2_120[14],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1934,addr_remain3_1934);


wire[15:0] addr_selector3_1935;
wire[15:0] addr_remain3_1935;
address_decode_4 decoder_3_1935 = address_decode_4(addr_selector2_120[15],addr_remain2_120[15:0],addr_remain2_120,addr_selector3_1935,addr_remain3_1935);


wire[15:0] addr_selector3_1936;
wire[15:0] addr_remain3_1936;
address_decode_4 decoder_3_1936 = address_decode_4(addr_selector2_121[0],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1936,addr_remain3_1936);


wire[15:0] addr_selector3_1937;
wire[15:0] addr_remain3_1937;
address_decode_4 decoder_3_1937 = address_decode_4(addr_selector2_121[1],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1937,addr_remain3_1937);


wire[15:0] addr_selector3_1938;
wire[15:0] addr_remain3_1938;
address_decode_4 decoder_3_1938 = address_decode_4(addr_selector2_121[2],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1938,addr_remain3_1938);


wire[15:0] addr_selector3_1939;
wire[15:0] addr_remain3_1939;
address_decode_4 decoder_3_1939 = address_decode_4(addr_selector2_121[3],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1939,addr_remain3_1939);


wire[15:0] addr_selector3_1940;
wire[15:0] addr_remain3_1940;
address_decode_4 decoder_3_1940 = address_decode_4(addr_selector2_121[4],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1940,addr_remain3_1940);


wire[15:0] addr_selector3_1941;
wire[15:0] addr_remain3_1941;
address_decode_4 decoder_3_1941 = address_decode_4(addr_selector2_121[5],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1941,addr_remain3_1941);


wire[15:0] addr_selector3_1942;
wire[15:0] addr_remain3_1942;
address_decode_4 decoder_3_1942 = address_decode_4(addr_selector2_121[6],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1942,addr_remain3_1942);


wire[15:0] addr_selector3_1943;
wire[15:0] addr_remain3_1943;
address_decode_4 decoder_3_1943 = address_decode_4(addr_selector2_121[7],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1943,addr_remain3_1943);


wire[15:0] addr_selector3_1944;
wire[15:0] addr_remain3_1944;
address_decode_4 decoder_3_1944 = address_decode_4(addr_selector2_121[8],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1944,addr_remain3_1944);


wire[15:0] addr_selector3_1945;
wire[15:0] addr_remain3_1945;
address_decode_4 decoder_3_1945 = address_decode_4(addr_selector2_121[9],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1945,addr_remain3_1945);


wire[15:0] addr_selector3_1946;
wire[15:0] addr_remain3_1946;
address_decode_4 decoder_3_1946 = address_decode_4(addr_selector2_121[10],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1946,addr_remain3_1946);


wire[15:0] addr_selector3_1947;
wire[15:0] addr_remain3_1947;
address_decode_4 decoder_3_1947 = address_decode_4(addr_selector2_121[11],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1947,addr_remain3_1947);


wire[15:0] addr_selector3_1948;
wire[15:0] addr_remain3_1948;
address_decode_4 decoder_3_1948 = address_decode_4(addr_selector2_121[12],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1948,addr_remain3_1948);


wire[15:0] addr_selector3_1949;
wire[15:0] addr_remain3_1949;
address_decode_4 decoder_3_1949 = address_decode_4(addr_selector2_121[13],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1949,addr_remain3_1949);


wire[15:0] addr_selector3_1950;
wire[15:0] addr_remain3_1950;
address_decode_4 decoder_3_1950 = address_decode_4(addr_selector2_121[14],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1950,addr_remain3_1950);


wire[15:0] addr_selector3_1951;
wire[15:0] addr_remain3_1951;
address_decode_4 decoder_3_1951 = address_decode_4(addr_selector2_121[15],addr_remain2_121[15:0],addr_remain2_121,addr_selector3_1951,addr_remain3_1951);


wire[15:0] addr_selector3_1952;
wire[15:0] addr_remain3_1952;
address_decode_4 decoder_3_1952 = address_decode_4(addr_selector2_122[0],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1952,addr_remain3_1952);


wire[15:0] addr_selector3_1953;
wire[15:0] addr_remain3_1953;
address_decode_4 decoder_3_1953 = address_decode_4(addr_selector2_122[1],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1953,addr_remain3_1953);


wire[15:0] addr_selector3_1954;
wire[15:0] addr_remain3_1954;
address_decode_4 decoder_3_1954 = address_decode_4(addr_selector2_122[2],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1954,addr_remain3_1954);


wire[15:0] addr_selector3_1955;
wire[15:0] addr_remain3_1955;
address_decode_4 decoder_3_1955 = address_decode_4(addr_selector2_122[3],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1955,addr_remain3_1955);


wire[15:0] addr_selector3_1956;
wire[15:0] addr_remain3_1956;
address_decode_4 decoder_3_1956 = address_decode_4(addr_selector2_122[4],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1956,addr_remain3_1956);


wire[15:0] addr_selector3_1957;
wire[15:0] addr_remain3_1957;
address_decode_4 decoder_3_1957 = address_decode_4(addr_selector2_122[5],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1957,addr_remain3_1957);


wire[15:0] addr_selector3_1958;
wire[15:0] addr_remain3_1958;
address_decode_4 decoder_3_1958 = address_decode_4(addr_selector2_122[6],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1958,addr_remain3_1958);


wire[15:0] addr_selector3_1959;
wire[15:0] addr_remain3_1959;
address_decode_4 decoder_3_1959 = address_decode_4(addr_selector2_122[7],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1959,addr_remain3_1959);


wire[15:0] addr_selector3_1960;
wire[15:0] addr_remain3_1960;
address_decode_4 decoder_3_1960 = address_decode_4(addr_selector2_122[8],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1960,addr_remain3_1960);


wire[15:0] addr_selector3_1961;
wire[15:0] addr_remain3_1961;
address_decode_4 decoder_3_1961 = address_decode_4(addr_selector2_122[9],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1961,addr_remain3_1961);


wire[15:0] addr_selector3_1962;
wire[15:0] addr_remain3_1962;
address_decode_4 decoder_3_1962 = address_decode_4(addr_selector2_122[10],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1962,addr_remain3_1962);


wire[15:0] addr_selector3_1963;
wire[15:0] addr_remain3_1963;
address_decode_4 decoder_3_1963 = address_decode_4(addr_selector2_122[11],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1963,addr_remain3_1963);


wire[15:0] addr_selector3_1964;
wire[15:0] addr_remain3_1964;
address_decode_4 decoder_3_1964 = address_decode_4(addr_selector2_122[12],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1964,addr_remain3_1964);


wire[15:0] addr_selector3_1965;
wire[15:0] addr_remain3_1965;
address_decode_4 decoder_3_1965 = address_decode_4(addr_selector2_122[13],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1965,addr_remain3_1965);


wire[15:0] addr_selector3_1966;
wire[15:0] addr_remain3_1966;
address_decode_4 decoder_3_1966 = address_decode_4(addr_selector2_122[14],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1966,addr_remain3_1966);


wire[15:0] addr_selector3_1967;
wire[15:0] addr_remain3_1967;
address_decode_4 decoder_3_1967 = address_decode_4(addr_selector2_122[15],addr_remain2_122[15:0],addr_remain2_122,addr_selector3_1967,addr_remain3_1967);


wire[15:0] addr_selector3_1968;
wire[15:0] addr_remain3_1968;
address_decode_4 decoder_3_1968 = address_decode_4(addr_selector2_123[0],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1968,addr_remain3_1968);


wire[15:0] addr_selector3_1969;
wire[15:0] addr_remain3_1969;
address_decode_4 decoder_3_1969 = address_decode_4(addr_selector2_123[1],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1969,addr_remain3_1969);


wire[15:0] addr_selector3_1970;
wire[15:0] addr_remain3_1970;
address_decode_4 decoder_3_1970 = address_decode_4(addr_selector2_123[2],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1970,addr_remain3_1970);


wire[15:0] addr_selector3_1971;
wire[15:0] addr_remain3_1971;
address_decode_4 decoder_3_1971 = address_decode_4(addr_selector2_123[3],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1971,addr_remain3_1971);


wire[15:0] addr_selector3_1972;
wire[15:0] addr_remain3_1972;
address_decode_4 decoder_3_1972 = address_decode_4(addr_selector2_123[4],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1972,addr_remain3_1972);


wire[15:0] addr_selector3_1973;
wire[15:0] addr_remain3_1973;
address_decode_4 decoder_3_1973 = address_decode_4(addr_selector2_123[5],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1973,addr_remain3_1973);


wire[15:0] addr_selector3_1974;
wire[15:0] addr_remain3_1974;
address_decode_4 decoder_3_1974 = address_decode_4(addr_selector2_123[6],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1974,addr_remain3_1974);


wire[15:0] addr_selector3_1975;
wire[15:0] addr_remain3_1975;
address_decode_4 decoder_3_1975 = address_decode_4(addr_selector2_123[7],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1975,addr_remain3_1975);


wire[15:0] addr_selector3_1976;
wire[15:0] addr_remain3_1976;
address_decode_4 decoder_3_1976 = address_decode_4(addr_selector2_123[8],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1976,addr_remain3_1976);


wire[15:0] addr_selector3_1977;
wire[15:0] addr_remain3_1977;
address_decode_4 decoder_3_1977 = address_decode_4(addr_selector2_123[9],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1977,addr_remain3_1977);


wire[15:0] addr_selector3_1978;
wire[15:0] addr_remain3_1978;
address_decode_4 decoder_3_1978 = address_decode_4(addr_selector2_123[10],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1978,addr_remain3_1978);


wire[15:0] addr_selector3_1979;
wire[15:0] addr_remain3_1979;
address_decode_4 decoder_3_1979 = address_decode_4(addr_selector2_123[11],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1979,addr_remain3_1979);


wire[15:0] addr_selector3_1980;
wire[15:0] addr_remain3_1980;
address_decode_4 decoder_3_1980 = address_decode_4(addr_selector2_123[12],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1980,addr_remain3_1980);


wire[15:0] addr_selector3_1981;
wire[15:0] addr_remain3_1981;
address_decode_4 decoder_3_1981 = address_decode_4(addr_selector2_123[13],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1981,addr_remain3_1981);


wire[15:0] addr_selector3_1982;
wire[15:0] addr_remain3_1982;
address_decode_4 decoder_3_1982 = address_decode_4(addr_selector2_123[14],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1982,addr_remain3_1982);


wire[15:0] addr_selector3_1983;
wire[15:0] addr_remain3_1983;
address_decode_4 decoder_3_1983 = address_decode_4(addr_selector2_123[15],addr_remain2_123[15:0],addr_remain2_123,addr_selector3_1983,addr_remain3_1983);


wire[15:0] addr_selector3_1984;
wire[15:0] addr_remain3_1984;
address_decode_4 decoder_3_1984 = address_decode_4(addr_selector2_124[0],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1984,addr_remain3_1984);


wire[15:0] addr_selector3_1985;
wire[15:0] addr_remain3_1985;
address_decode_4 decoder_3_1985 = address_decode_4(addr_selector2_124[1],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1985,addr_remain3_1985);


wire[15:0] addr_selector3_1986;
wire[15:0] addr_remain3_1986;
address_decode_4 decoder_3_1986 = address_decode_4(addr_selector2_124[2],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1986,addr_remain3_1986);


wire[15:0] addr_selector3_1987;
wire[15:0] addr_remain3_1987;
address_decode_4 decoder_3_1987 = address_decode_4(addr_selector2_124[3],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1987,addr_remain3_1987);


wire[15:0] addr_selector3_1988;
wire[15:0] addr_remain3_1988;
address_decode_4 decoder_3_1988 = address_decode_4(addr_selector2_124[4],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1988,addr_remain3_1988);


wire[15:0] addr_selector3_1989;
wire[15:0] addr_remain3_1989;
address_decode_4 decoder_3_1989 = address_decode_4(addr_selector2_124[5],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1989,addr_remain3_1989);


wire[15:0] addr_selector3_1990;
wire[15:0] addr_remain3_1990;
address_decode_4 decoder_3_1990 = address_decode_4(addr_selector2_124[6],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1990,addr_remain3_1990);


wire[15:0] addr_selector3_1991;
wire[15:0] addr_remain3_1991;
address_decode_4 decoder_3_1991 = address_decode_4(addr_selector2_124[7],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1991,addr_remain3_1991);


wire[15:0] addr_selector3_1992;
wire[15:0] addr_remain3_1992;
address_decode_4 decoder_3_1992 = address_decode_4(addr_selector2_124[8],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1992,addr_remain3_1992);


wire[15:0] addr_selector3_1993;
wire[15:0] addr_remain3_1993;
address_decode_4 decoder_3_1993 = address_decode_4(addr_selector2_124[9],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1993,addr_remain3_1993);


wire[15:0] addr_selector3_1994;
wire[15:0] addr_remain3_1994;
address_decode_4 decoder_3_1994 = address_decode_4(addr_selector2_124[10],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1994,addr_remain3_1994);


wire[15:0] addr_selector3_1995;
wire[15:0] addr_remain3_1995;
address_decode_4 decoder_3_1995 = address_decode_4(addr_selector2_124[11],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1995,addr_remain3_1995);


wire[15:0] addr_selector3_1996;
wire[15:0] addr_remain3_1996;
address_decode_4 decoder_3_1996 = address_decode_4(addr_selector2_124[12],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1996,addr_remain3_1996);


wire[15:0] addr_selector3_1997;
wire[15:0] addr_remain3_1997;
address_decode_4 decoder_3_1997 = address_decode_4(addr_selector2_124[13],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1997,addr_remain3_1997);


wire[15:0] addr_selector3_1998;
wire[15:0] addr_remain3_1998;
address_decode_4 decoder_3_1998 = address_decode_4(addr_selector2_124[14],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1998,addr_remain3_1998);


wire[15:0] addr_selector3_1999;
wire[15:0] addr_remain3_1999;
address_decode_4 decoder_3_1999 = address_decode_4(addr_selector2_124[15],addr_remain2_124[15:0],addr_remain2_124,addr_selector3_1999,addr_remain3_1999);


wire[15:0] addr_selector3_2000;
wire[15:0] addr_remain3_2000;
address_decode_4 decoder_3_2000 = address_decode_4(addr_selector2_125[0],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2000,addr_remain3_2000);


wire[15:0] addr_selector3_2001;
wire[15:0] addr_remain3_2001;
address_decode_4 decoder_3_2001 = address_decode_4(addr_selector2_125[1],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2001,addr_remain3_2001);


wire[15:0] addr_selector3_2002;
wire[15:0] addr_remain3_2002;
address_decode_4 decoder_3_2002 = address_decode_4(addr_selector2_125[2],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2002,addr_remain3_2002);


wire[15:0] addr_selector3_2003;
wire[15:0] addr_remain3_2003;
address_decode_4 decoder_3_2003 = address_decode_4(addr_selector2_125[3],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2003,addr_remain3_2003);


wire[15:0] addr_selector3_2004;
wire[15:0] addr_remain3_2004;
address_decode_4 decoder_3_2004 = address_decode_4(addr_selector2_125[4],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2004,addr_remain3_2004);


wire[15:0] addr_selector3_2005;
wire[15:0] addr_remain3_2005;
address_decode_4 decoder_3_2005 = address_decode_4(addr_selector2_125[5],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2005,addr_remain3_2005);


wire[15:0] addr_selector3_2006;
wire[15:0] addr_remain3_2006;
address_decode_4 decoder_3_2006 = address_decode_4(addr_selector2_125[6],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2006,addr_remain3_2006);


wire[15:0] addr_selector3_2007;
wire[15:0] addr_remain3_2007;
address_decode_4 decoder_3_2007 = address_decode_4(addr_selector2_125[7],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2007,addr_remain3_2007);


wire[15:0] addr_selector3_2008;
wire[15:0] addr_remain3_2008;
address_decode_4 decoder_3_2008 = address_decode_4(addr_selector2_125[8],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2008,addr_remain3_2008);


wire[15:0] addr_selector3_2009;
wire[15:0] addr_remain3_2009;
address_decode_4 decoder_3_2009 = address_decode_4(addr_selector2_125[9],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2009,addr_remain3_2009);


wire[15:0] addr_selector3_2010;
wire[15:0] addr_remain3_2010;
address_decode_4 decoder_3_2010 = address_decode_4(addr_selector2_125[10],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2010,addr_remain3_2010);


wire[15:0] addr_selector3_2011;
wire[15:0] addr_remain3_2011;
address_decode_4 decoder_3_2011 = address_decode_4(addr_selector2_125[11],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2011,addr_remain3_2011);


wire[15:0] addr_selector3_2012;
wire[15:0] addr_remain3_2012;
address_decode_4 decoder_3_2012 = address_decode_4(addr_selector2_125[12],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2012,addr_remain3_2012);


wire[15:0] addr_selector3_2013;
wire[15:0] addr_remain3_2013;
address_decode_4 decoder_3_2013 = address_decode_4(addr_selector2_125[13],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2013,addr_remain3_2013);


wire[15:0] addr_selector3_2014;
wire[15:0] addr_remain3_2014;
address_decode_4 decoder_3_2014 = address_decode_4(addr_selector2_125[14],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2014,addr_remain3_2014);


wire[15:0] addr_selector3_2015;
wire[15:0] addr_remain3_2015;
address_decode_4 decoder_3_2015 = address_decode_4(addr_selector2_125[15],addr_remain2_125[15:0],addr_remain2_125,addr_selector3_2015,addr_remain3_2015);


wire[15:0] addr_selector3_2016;
wire[15:0] addr_remain3_2016;
address_decode_4 decoder_3_2016 = address_decode_4(addr_selector2_126[0],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2016,addr_remain3_2016);


wire[15:0] addr_selector3_2017;
wire[15:0] addr_remain3_2017;
address_decode_4 decoder_3_2017 = address_decode_4(addr_selector2_126[1],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2017,addr_remain3_2017);


wire[15:0] addr_selector3_2018;
wire[15:0] addr_remain3_2018;
address_decode_4 decoder_3_2018 = address_decode_4(addr_selector2_126[2],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2018,addr_remain3_2018);


wire[15:0] addr_selector3_2019;
wire[15:0] addr_remain3_2019;
address_decode_4 decoder_3_2019 = address_decode_4(addr_selector2_126[3],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2019,addr_remain3_2019);


wire[15:0] addr_selector3_2020;
wire[15:0] addr_remain3_2020;
address_decode_4 decoder_3_2020 = address_decode_4(addr_selector2_126[4],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2020,addr_remain3_2020);


wire[15:0] addr_selector3_2021;
wire[15:0] addr_remain3_2021;
address_decode_4 decoder_3_2021 = address_decode_4(addr_selector2_126[5],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2021,addr_remain3_2021);


wire[15:0] addr_selector3_2022;
wire[15:0] addr_remain3_2022;
address_decode_4 decoder_3_2022 = address_decode_4(addr_selector2_126[6],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2022,addr_remain3_2022);


wire[15:0] addr_selector3_2023;
wire[15:0] addr_remain3_2023;
address_decode_4 decoder_3_2023 = address_decode_4(addr_selector2_126[7],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2023,addr_remain3_2023);


wire[15:0] addr_selector3_2024;
wire[15:0] addr_remain3_2024;
address_decode_4 decoder_3_2024 = address_decode_4(addr_selector2_126[8],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2024,addr_remain3_2024);


wire[15:0] addr_selector3_2025;
wire[15:0] addr_remain3_2025;
address_decode_4 decoder_3_2025 = address_decode_4(addr_selector2_126[9],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2025,addr_remain3_2025);


wire[15:0] addr_selector3_2026;
wire[15:0] addr_remain3_2026;
address_decode_4 decoder_3_2026 = address_decode_4(addr_selector2_126[10],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2026,addr_remain3_2026);


wire[15:0] addr_selector3_2027;
wire[15:0] addr_remain3_2027;
address_decode_4 decoder_3_2027 = address_decode_4(addr_selector2_126[11],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2027,addr_remain3_2027);


wire[15:0] addr_selector3_2028;
wire[15:0] addr_remain3_2028;
address_decode_4 decoder_3_2028 = address_decode_4(addr_selector2_126[12],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2028,addr_remain3_2028);


wire[15:0] addr_selector3_2029;
wire[15:0] addr_remain3_2029;
address_decode_4 decoder_3_2029 = address_decode_4(addr_selector2_126[13],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2029,addr_remain3_2029);


wire[15:0] addr_selector3_2030;
wire[15:0] addr_remain3_2030;
address_decode_4 decoder_3_2030 = address_decode_4(addr_selector2_126[14],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2030,addr_remain3_2030);


wire[15:0] addr_selector3_2031;
wire[15:0] addr_remain3_2031;
address_decode_4 decoder_3_2031 = address_decode_4(addr_selector2_126[15],addr_remain2_126[15:0],addr_remain2_126,addr_selector3_2031,addr_remain3_2031);


wire[15:0] addr_selector3_2032;
wire[15:0] addr_remain3_2032;
address_decode_4 decoder_3_2032 = address_decode_4(addr_selector2_127[0],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2032,addr_remain3_2032);


wire[15:0] addr_selector3_2033;
wire[15:0] addr_remain3_2033;
address_decode_4 decoder_3_2033 = address_decode_4(addr_selector2_127[1],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2033,addr_remain3_2033);


wire[15:0] addr_selector3_2034;
wire[15:0] addr_remain3_2034;
address_decode_4 decoder_3_2034 = address_decode_4(addr_selector2_127[2],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2034,addr_remain3_2034);


wire[15:0] addr_selector3_2035;
wire[15:0] addr_remain3_2035;
address_decode_4 decoder_3_2035 = address_decode_4(addr_selector2_127[3],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2035,addr_remain3_2035);


wire[15:0] addr_selector3_2036;
wire[15:0] addr_remain3_2036;
address_decode_4 decoder_3_2036 = address_decode_4(addr_selector2_127[4],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2036,addr_remain3_2036);


wire[15:0] addr_selector3_2037;
wire[15:0] addr_remain3_2037;
address_decode_4 decoder_3_2037 = address_decode_4(addr_selector2_127[5],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2037,addr_remain3_2037);


wire[15:0] addr_selector3_2038;
wire[15:0] addr_remain3_2038;
address_decode_4 decoder_3_2038 = address_decode_4(addr_selector2_127[6],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2038,addr_remain3_2038);


wire[15:0] addr_selector3_2039;
wire[15:0] addr_remain3_2039;
address_decode_4 decoder_3_2039 = address_decode_4(addr_selector2_127[7],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2039,addr_remain3_2039);


wire[15:0] addr_selector3_2040;
wire[15:0] addr_remain3_2040;
address_decode_4 decoder_3_2040 = address_decode_4(addr_selector2_127[8],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2040,addr_remain3_2040);


wire[15:0] addr_selector3_2041;
wire[15:0] addr_remain3_2041;
address_decode_4 decoder_3_2041 = address_decode_4(addr_selector2_127[9],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2041,addr_remain3_2041);


wire[15:0] addr_selector3_2042;
wire[15:0] addr_remain3_2042;
address_decode_4 decoder_3_2042 = address_decode_4(addr_selector2_127[10],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2042,addr_remain3_2042);


wire[15:0] addr_selector3_2043;
wire[15:0] addr_remain3_2043;
address_decode_4 decoder_3_2043 = address_decode_4(addr_selector2_127[11],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2043,addr_remain3_2043);


wire[15:0] addr_selector3_2044;
wire[15:0] addr_remain3_2044;
address_decode_4 decoder_3_2044 = address_decode_4(addr_selector2_127[12],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2044,addr_remain3_2044);


wire[15:0] addr_selector3_2045;
wire[15:0] addr_remain3_2045;
address_decode_4 decoder_3_2045 = address_decode_4(addr_selector2_127[13],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2045,addr_remain3_2045);


wire[15:0] addr_selector3_2046;
wire[15:0] addr_remain3_2046;
address_decode_4 decoder_3_2046 = address_decode_4(addr_selector2_127[14],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2046,addr_remain3_2046);


wire[15:0] addr_selector3_2047;
wire[15:0] addr_remain3_2047;
address_decode_4 decoder_3_2047 = address_decode_4(addr_selector2_127[15],addr_remain2_127[15:0],addr_remain2_127,addr_selector3_2047,addr_remain3_2047);


wire[15:0] addr_selector3_2048;
wire[15:0] addr_remain3_2048;
address_decode_4 decoder_3_2048 = address_decode_4(addr_selector2_128[0],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2048,addr_remain3_2048);


wire[15:0] addr_selector3_2049;
wire[15:0] addr_remain3_2049;
address_decode_4 decoder_3_2049 = address_decode_4(addr_selector2_128[1],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2049,addr_remain3_2049);


wire[15:0] addr_selector3_2050;
wire[15:0] addr_remain3_2050;
address_decode_4 decoder_3_2050 = address_decode_4(addr_selector2_128[2],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2050,addr_remain3_2050);


wire[15:0] addr_selector3_2051;
wire[15:0] addr_remain3_2051;
address_decode_4 decoder_3_2051 = address_decode_4(addr_selector2_128[3],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2051,addr_remain3_2051);


wire[15:0] addr_selector3_2052;
wire[15:0] addr_remain3_2052;
address_decode_4 decoder_3_2052 = address_decode_4(addr_selector2_128[4],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2052,addr_remain3_2052);


wire[15:0] addr_selector3_2053;
wire[15:0] addr_remain3_2053;
address_decode_4 decoder_3_2053 = address_decode_4(addr_selector2_128[5],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2053,addr_remain3_2053);


wire[15:0] addr_selector3_2054;
wire[15:0] addr_remain3_2054;
address_decode_4 decoder_3_2054 = address_decode_4(addr_selector2_128[6],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2054,addr_remain3_2054);


wire[15:0] addr_selector3_2055;
wire[15:0] addr_remain3_2055;
address_decode_4 decoder_3_2055 = address_decode_4(addr_selector2_128[7],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2055,addr_remain3_2055);


wire[15:0] addr_selector3_2056;
wire[15:0] addr_remain3_2056;
address_decode_4 decoder_3_2056 = address_decode_4(addr_selector2_128[8],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2056,addr_remain3_2056);


wire[15:0] addr_selector3_2057;
wire[15:0] addr_remain3_2057;
address_decode_4 decoder_3_2057 = address_decode_4(addr_selector2_128[9],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2057,addr_remain3_2057);


wire[15:0] addr_selector3_2058;
wire[15:0] addr_remain3_2058;
address_decode_4 decoder_3_2058 = address_decode_4(addr_selector2_128[10],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2058,addr_remain3_2058);


wire[15:0] addr_selector3_2059;
wire[15:0] addr_remain3_2059;
address_decode_4 decoder_3_2059 = address_decode_4(addr_selector2_128[11],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2059,addr_remain3_2059);


wire[15:0] addr_selector3_2060;
wire[15:0] addr_remain3_2060;
address_decode_4 decoder_3_2060 = address_decode_4(addr_selector2_128[12],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2060,addr_remain3_2060);


wire[15:0] addr_selector3_2061;
wire[15:0] addr_remain3_2061;
address_decode_4 decoder_3_2061 = address_decode_4(addr_selector2_128[13],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2061,addr_remain3_2061);


wire[15:0] addr_selector3_2062;
wire[15:0] addr_remain3_2062;
address_decode_4 decoder_3_2062 = address_decode_4(addr_selector2_128[14],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2062,addr_remain3_2062);


wire[15:0] addr_selector3_2063;
wire[15:0] addr_remain3_2063;
address_decode_4 decoder_3_2063 = address_decode_4(addr_selector2_128[15],addr_remain2_128[15:0],addr_remain2_128,addr_selector3_2063,addr_remain3_2063);


wire[15:0] addr_selector3_2064;
wire[15:0] addr_remain3_2064;
address_decode_4 decoder_3_2064 = address_decode_4(addr_selector2_129[0],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2064,addr_remain3_2064);


wire[15:0] addr_selector3_2065;
wire[15:0] addr_remain3_2065;
address_decode_4 decoder_3_2065 = address_decode_4(addr_selector2_129[1],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2065,addr_remain3_2065);


wire[15:0] addr_selector3_2066;
wire[15:0] addr_remain3_2066;
address_decode_4 decoder_3_2066 = address_decode_4(addr_selector2_129[2],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2066,addr_remain3_2066);


wire[15:0] addr_selector3_2067;
wire[15:0] addr_remain3_2067;
address_decode_4 decoder_3_2067 = address_decode_4(addr_selector2_129[3],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2067,addr_remain3_2067);


wire[15:0] addr_selector3_2068;
wire[15:0] addr_remain3_2068;
address_decode_4 decoder_3_2068 = address_decode_4(addr_selector2_129[4],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2068,addr_remain3_2068);


wire[15:0] addr_selector3_2069;
wire[15:0] addr_remain3_2069;
address_decode_4 decoder_3_2069 = address_decode_4(addr_selector2_129[5],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2069,addr_remain3_2069);


wire[15:0] addr_selector3_2070;
wire[15:0] addr_remain3_2070;
address_decode_4 decoder_3_2070 = address_decode_4(addr_selector2_129[6],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2070,addr_remain3_2070);


wire[15:0] addr_selector3_2071;
wire[15:0] addr_remain3_2071;
address_decode_4 decoder_3_2071 = address_decode_4(addr_selector2_129[7],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2071,addr_remain3_2071);


wire[15:0] addr_selector3_2072;
wire[15:0] addr_remain3_2072;
address_decode_4 decoder_3_2072 = address_decode_4(addr_selector2_129[8],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2072,addr_remain3_2072);


wire[15:0] addr_selector3_2073;
wire[15:0] addr_remain3_2073;
address_decode_4 decoder_3_2073 = address_decode_4(addr_selector2_129[9],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2073,addr_remain3_2073);


wire[15:0] addr_selector3_2074;
wire[15:0] addr_remain3_2074;
address_decode_4 decoder_3_2074 = address_decode_4(addr_selector2_129[10],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2074,addr_remain3_2074);


wire[15:0] addr_selector3_2075;
wire[15:0] addr_remain3_2075;
address_decode_4 decoder_3_2075 = address_decode_4(addr_selector2_129[11],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2075,addr_remain3_2075);


wire[15:0] addr_selector3_2076;
wire[15:0] addr_remain3_2076;
address_decode_4 decoder_3_2076 = address_decode_4(addr_selector2_129[12],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2076,addr_remain3_2076);


wire[15:0] addr_selector3_2077;
wire[15:0] addr_remain3_2077;
address_decode_4 decoder_3_2077 = address_decode_4(addr_selector2_129[13],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2077,addr_remain3_2077);


wire[15:0] addr_selector3_2078;
wire[15:0] addr_remain3_2078;
address_decode_4 decoder_3_2078 = address_decode_4(addr_selector2_129[14],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2078,addr_remain3_2078);


wire[15:0] addr_selector3_2079;
wire[15:0] addr_remain3_2079;
address_decode_4 decoder_3_2079 = address_decode_4(addr_selector2_129[15],addr_remain2_129[15:0],addr_remain2_129,addr_selector3_2079,addr_remain3_2079);


wire[15:0] addr_selector3_2080;
wire[15:0] addr_remain3_2080;
address_decode_4 decoder_3_2080 = address_decode_4(addr_selector2_130[0],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2080,addr_remain3_2080);


wire[15:0] addr_selector3_2081;
wire[15:0] addr_remain3_2081;
address_decode_4 decoder_3_2081 = address_decode_4(addr_selector2_130[1],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2081,addr_remain3_2081);


wire[15:0] addr_selector3_2082;
wire[15:0] addr_remain3_2082;
address_decode_4 decoder_3_2082 = address_decode_4(addr_selector2_130[2],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2082,addr_remain3_2082);


wire[15:0] addr_selector3_2083;
wire[15:0] addr_remain3_2083;
address_decode_4 decoder_3_2083 = address_decode_4(addr_selector2_130[3],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2083,addr_remain3_2083);


wire[15:0] addr_selector3_2084;
wire[15:0] addr_remain3_2084;
address_decode_4 decoder_3_2084 = address_decode_4(addr_selector2_130[4],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2084,addr_remain3_2084);


wire[15:0] addr_selector3_2085;
wire[15:0] addr_remain3_2085;
address_decode_4 decoder_3_2085 = address_decode_4(addr_selector2_130[5],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2085,addr_remain3_2085);


wire[15:0] addr_selector3_2086;
wire[15:0] addr_remain3_2086;
address_decode_4 decoder_3_2086 = address_decode_4(addr_selector2_130[6],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2086,addr_remain3_2086);


wire[15:0] addr_selector3_2087;
wire[15:0] addr_remain3_2087;
address_decode_4 decoder_3_2087 = address_decode_4(addr_selector2_130[7],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2087,addr_remain3_2087);


wire[15:0] addr_selector3_2088;
wire[15:0] addr_remain3_2088;
address_decode_4 decoder_3_2088 = address_decode_4(addr_selector2_130[8],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2088,addr_remain3_2088);


wire[15:0] addr_selector3_2089;
wire[15:0] addr_remain3_2089;
address_decode_4 decoder_3_2089 = address_decode_4(addr_selector2_130[9],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2089,addr_remain3_2089);


wire[15:0] addr_selector3_2090;
wire[15:0] addr_remain3_2090;
address_decode_4 decoder_3_2090 = address_decode_4(addr_selector2_130[10],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2090,addr_remain3_2090);


wire[15:0] addr_selector3_2091;
wire[15:0] addr_remain3_2091;
address_decode_4 decoder_3_2091 = address_decode_4(addr_selector2_130[11],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2091,addr_remain3_2091);


wire[15:0] addr_selector3_2092;
wire[15:0] addr_remain3_2092;
address_decode_4 decoder_3_2092 = address_decode_4(addr_selector2_130[12],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2092,addr_remain3_2092);


wire[15:0] addr_selector3_2093;
wire[15:0] addr_remain3_2093;
address_decode_4 decoder_3_2093 = address_decode_4(addr_selector2_130[13],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2093,addr_remain3_2093);


wire[15:0] addr_selector3_2094;
wire[15:0] addr_remain3_2094;
address_decode_4 decoder_3_2094 = address_decode_4(addr_selector2_130[14],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2094,addr_remain3_2094);


wire[15:0] addr_selector3_2095;
wire[15:0] addr_remain3_2095;
address_decode_4 decoder_3_2095 = address_decode_4(addr_selector2_130[15],addr_remain2_130[15:0],addr_remain2_130,addr_selector3_2095,addr_remain3_2095);


wire[15:0] addr_selector3_2096;
wire[15:0] addr_remain3_2096;
address_decode_4 decoder_3_2096 = address_decode_4(addr_selector2_131[0],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2096,addr_remain3_2096);


wire[15:0] addr_selector3_2097;
wire[15:0] addr_remain3_2097;
address_decode_4 decoder_3_2097 = address_decode_4(addr_selector2_131[1],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2097,addr_remain3_2097);


wire[15:0] addr_selector3_2098;
wire[15:0] addr_remain3_2098;
address_decode_4 decoder_3_2098 = address_decode_4(addr_selector2_131[2],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2098,addr_remain3_2098);


wire[15:0] addr_selector3_2099;
wire[15:0] addr_remain3_2099;
address_decode_4 decoder_3_2099 = address_decode_4(addr_selector2_131[3],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2099,addr_remain3_2099);


wire[15:0] addr_selector3_2100;
wire[15:0] addr_remain3_2100;
address_decode_4 decoder_3_2100 = address_decode_4(addr_selector2_131[4],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2100,addr_remain3_2100);


wire[15:0] addr_selector3_2101;
wire[15:0] addr_remain3_2101;
address_decode_4 decoder_3_2101 = address_decode_4(addr_selector2_131[5],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2101,addr_remain3_2101);


wire[15:0] addr_selector3_2102;
wire[15:0] addr_remain3_2102;
address_decode_4 decoder_3_2102 = address_decode_4(addr_selector2_131[6],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2102,addr_remain3_2102);


wire[15:0] addr_selector3_2103;
wire[15:0] addr_remain3_2103;
address_decode_4 decoder_3_2103 = address_decode_4(addr_selector2_131[7],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2103,addr_remain3_2103);


wire[15:0] addr_selector3_2104;
wire[15:0] addr_remain3_2104;
address_decode_4 decoder_3_2104 = address_decode_4(addr_selector2_131[8],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2104,addr_remain3_2104);


wire[15:0] addr_selector3_2105;
wire[15:0] addr_remain3_2105;
address_decode_4 decoder_3_2105 = address_decode_4(addr_selector2_131[9],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2105,addr_remain3_2105);


wire[15:0] addr_selector3_2106;
wire[15:0] addr_remain3_2106;
address_decode_4 decoder_3_2106 = address_decode_4(addr_selector2_131[10],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2106,addr_remain3_2106);


wire[15:0] addr_selector3_2107;
wire[15:0] addr_remain3_2107;
address_decode_4 decoder_3_2107 = address_decode_4(addr_selector2_131[11],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2107,addr_remain3_2107);


wire[15:0] addr_selector3_2108;
wire[15:0] addr_remain3_2108;
address_decode_4 decoder_3_2108 = address_decode_4(addr_selector2_131[12],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2108,addr_remain3_2108);


wire[15:0] addr_selector3_2109;
wire[15:0] addr_remain3_2109;
address_decode_4 decoder_3_2109 = address_decode_4(addr_selector2_131[13],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2109,addr_remain3_2109);


wire[15:0] addr_selector3_2110;
wire[15:0] addr_remain3_2110;
address_decode_4 decoder_3_2110 = address_decode_4(addr_selector2_131[14],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2110,addr_remain3_2110);


wire[15:0] addr_selector3_2111;
wire[15:0] addr_remain3_2111;
address_decode_4 decoder_3_2111 = address_decode_4(addr_selector2_131[15],addr_remain2_131[15:0],addr_remain2_131,addr_selector3_2111,addr_remain3_2111);


wire[15:0] addr_selector3_2112;
wire[15:0] addr_remain3_2112;
address_decode_4 decoder_3_2112 = address_decode_4(addr_selector2_132[0],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2112,addr_remain3_2112);


wire[15:0] addr_selector3_2113;
wire[15:0] addr_remain3_2113;
address_decode_4 decoder_3_2113 = address_decode_4(addr_selector2_132[1],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2113,addr_remain3_2113);


wire[15:0] addr_selector3_2114;
wire[15:0] addr_remain3_2114;
address_decode_4 decoder_3_2114 = address_decode_4(addr_selector2_132[2],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2114,addr_remain3_2114);


wire[15:0] addr_selector3_2115;
wire[15:0] addr_remain3_2115;
address_decode_4 decoder_3_2115 = address_decode_4(addr_selector2_132[3],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2115,addr_remain3_2115);


wire[15:0] addr_selector3_2116;
wire[15:0] addr_remain3_2116;
address_decode_4 decoder_3_2116 = address_decode_4(addr_selector2_132[4],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2116,addr_remain3_2116);


wire[15:0] addr_selector3_2117;
wire[15:0] addr_remain3_2117;
address_decode_4 decoder_3_2117 = address_decode_4(addr_selector2_132[5],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2117,addr_remain3_2117);


wire[15:0] addr_selector3_2118;
wire[15:0] addr_remain3_2118;
address_decode_4 decoder_3_2118 = address_decode_4(addr_selector2_132[6],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2118,addr_remain3_2118);


wire[15:0] addr_selector3_2119;
wire[15:0] addr_remain3_2119;
address_decode_4 decoder_3_2119 = address_decode_4(addr_selector2_132[7],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2119,addr_remain3_2119);


wire[15:0] addr_selector3_2120;
wire[15:0] addr_remain3_2120;
address_decode_4 decoder_3_2120 = address_decode_4(addr_selector2_132[8],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2120,addr_remain3_2120);


wire[15:0] addr_selector3_2121;
wire[15:0] addr_remain3_2121;
address_decode_4 decoder_3_2121 = address_decode_4(addr_selector2_132[9],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2121,addr_remain3_2121);


wire[15:0] addr_selector3_2122;
wire[15:0] addr_remain3_2122;
address_decode_4 decoder_3_2122 = address_decode_4(addr_selector2_132[10],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2122,addr_remain3_2122);


wire[15:0] addr_selector3_2123;
wire[15:0] addr_remain3_2123;
address_decode_4 decoder_3_2123 = address_decode_4(addr_selector2_132[11],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2123,addr_remain3_2123);


wire[15:0] addr_selector3_2124;
wire[15:0] addr_remain3_2124;
address_decode_4 decoder_3_2124 = address_decode_4(addr_selector2_132[12],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2124,addr_remain3_2124);


wire[15:0] addr_selector3_2125;
wire[15:0] addr_remain3_2125;
address_decode_4 decoder_3_2125 = address_decode_4(addr_selector2_132[13],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2125,addr_remain3_2125);


wire[15:0] addr_selector3_2126;
wire[15:0] addr_remain3_2126;
address_decode_4 decoder_3_2126 = address_decode_4(addr_selector2_132[14],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2126,addr_remain3_2126);


wire[15:0] addr_selector3_2127;
wire[15:0] addr_remain3_2127;
address_decode_4 decoder_3_2127 = address_decode_4(addr_selector2_132[15],addr_remain2_132[15:0],addr_remain2_132,addr_selector3_2127,addr_remain3_2127);


wire[15:0] addr_selector3_2128;
wire[15:0] addr_remain3_2128;
address_decode_4 decoder_3_2128 = address_decode_4(addr_selector2_133[0],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2128,addr_remain3_2128);


wire[15:0] addr_selector3_2129;
wire[15:0] addr_remain3_2129;
address_decode_4 decoder_3_2129 = address_decode_4(addr_selector2_133[1],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2129,addr_remain3_2129);


wire[15:0] addr_selector3_2130;
wire[15:0] addr_remain3_2130;
address_decode_4 decoder_3_2130 = address_decode_4(addr_selector2_133[2],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2130,addr_remain3_2130);


wire[15:0] addr_selector3_2131;
wire[15:0] addr_remain3_2131;
address_decode_4 decoder_3_2131 = address_decode_4(addr_selector2_133[3],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2131,addr_remain3_2131);


wire[15:0] addr_selector3_2132;
wire[15:0] addr_remain3_2132;
address_decode_4 decoder_3_2132 = address_decode_4(addr_selector2_133[4],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2132,addr_remain3_2132);


wire[15:0] addr_selector3_2133;
wire[15:0] addr_remain3_2133;
address_decode_4 decoder_3_2133 = address_decode_4(addr_selector2_133[5],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2133,addr_remain3_2133);


wire[15:0] addr_selector3_2134;
wire[15:0] addr_remain3_2134;
address_decode_4 decoder_3_2134 = address_decode_4(addr_selector2_133[6],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2134,addr_remain3_2134);


wire[15:0] addr_selector3_2135;
wire[15:0] addr_remain3_2135;
address_decode_4 decoder_3_2135 = address_decode_4(addr_selector2_133[7],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2135,addr_remain3_2135);


wire[15:0] addr_selector3_2136;
wire[15:0] addr_remain3_2136;
address_decode_4 decoder_3_2136 = address_decode_4(addr_selector2_133[8],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2136,addr_remain3_2136);


wire[15:0] addr_selector3_2137;
wire[15:0] addr_remain3_2137;
address_decode_4 decoder_3_2137 = address_decode_4(addr_selector2_133[9],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2137,addr_remain3_2137);


wire[15:0] addr_selector3_2138;
wire[15:0] addr_remain3_2138;
address_decode_4 decoder_3_2138 = address_decode_4(addr_selector2_133[10],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2138,addr_remain3_2138);


wire[15:0] addr_selector3_2139;
wire[15:0] addr_remain3_2139;
address_decode_4 decoder_3_2139 = address_decode_4(addr_selector2_133[11],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2139,addr_remain3_2139);


wire[15:0] addr_selector3_2140;
wire[15:0] addr_remain3_2140;
address_decode_4 decoder_3_2140 = address_decode_4(addr_selector2_133[12],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2140,addr_remain3_2140);


wire[15:0] addr_selector3_2141;
wire[15:0] addr_remain3_2141;
address_decode_4 decoder_3_2141 = address_decode_4(addr_selector2_133[13],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2141,addr_remain3_2141);


wire[15:0] addr_selector3_2142;
wire[15:0] addr_remain3_2142;
address_decode_4 decoder_3_2142 = address_decode_4(addr_selector2_133[14],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2142,addr_remain3_2142);


wire[15:0] addr_selector3_2143;
wire[15:0] addr_remain3_2143;
address_decode_4 decoder_3_2143 = address_decode_4(addr_selector2_133[15],addr_remain2_133[15:0],addr_remain2_133,addr_selector3_2143,addr_remain3_2143);


wire[15:0] addr_selector3_2144;
wire[15:0] addr_remain3_2144;
address_decode_4 decoder_3_2144 = address_decode_4(addr_selector2_134[0],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2144,addr_remain3_2144);


wire[15:0] addr_selector3_2145;
wire[15:0] addr_remain3_2145;
address_decode_4 decoder_3_2145 = address_decode_4(addr_selector2_134[1],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2145,addr_remain3_2145);


wire[15:0] addr_selector3_2146;
wire[15:0] addr_remain3_2146;
address_decode_4 decoder_3_2146 = address_decode_4(addr_selector2_134[2],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2146,addr_remain3_2146);


wire[15:0] addr_selector3_2147;
wire[15:0] addr_remain3_2147;
address_decode_4 decoder_3_2147 = address_decode_4(addr_selector2_134[3],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2147,addr_remain3_2147);


wire[15:0] addr_selector3_2148;
wire[15:0] addr_remain3_2148;
address_decode_4 decoder_3_2148 = address_decode_4(addr_selector2_134[4],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2148,addr_remain3_2148);


wire[15:0] addr_selector3_2149;
wire[15:0] addr_remain3_2149;
address_decode_4 decoder_3_2149 = address_decode_4(addr_selector2_134[5],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2149,addr_remain3_2149);


wire[15:0] addr_selector3_2150;
wire[15:0] addr_remain3_2150;
address_decode_4 decoder_3_2150 = address_decode_4(addr_selector2_134[6],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2150,addr_remain3_2150);


wire[15:0] addr_selector3_2151;
wire[15:0] addr_remain3_2151;
address_decode_4 decoder_3_2151 = address_decode_4(addr_selector2_134[7],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2151,addr_remain3_2151);


wire[15:0] addr_selector3_2152;
wire[15:0] addr_remain3_2152;
address_decode_4 decoder_3_2152 = address_decode_4(addr_selector2_134[8],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2152,addr_remain3_2152);


wire[15:0] addr_selector3_2153;
wire[15:0] addr_remain3_2153;
address_decode_4 decoder_3_2153 = address_decode_4(addr_selector2_134[9],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2153,addr_remain3_2153);


wire[15:0] addr_selector3_2154;
wire[15:0] addr_remain3_2154;
address_decode_4 decoder_3_2154 = address_decode_4(addr_selector2_134[10],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2154,addr_remain3_2154);


wire[15:0] addr_selector3_2155;
wire[15:0] addr_remain3_2155;
address_decode_4 decoder_3_2155 = address_decode_4(addr_selector2_134[11],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2155,addr_remain3_2155);


wire[15:0] addr_selector3_2156;
wire[15:0] addr_remain3_2156;
address_decode_4 decoder_3_2156 = address_decode_4(addr_selector2_134[12],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2156,addr_remain3_2156);


wire[15:0] addr_selector3_2157;
wire[15:0] addr_remain3_2157;
address_decode_4 decoder_3_2157 = address_decode_4(addr_selector2_134[13],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2157,addr_remain3_2157);


wire[15:0] addr_selector3_2158;
wire[15:0] addr_remain3_2158;
address_decode_4 decoder_3_2158 = address_decode_4(addr_selector2_134[14],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2158,addr_remain3_2158);


wire[15:0] addr_selector3_2159;
wire[15:0] addr_remain3_2159;
address_decode_4 decoder_3_2159 = address_decode_4(addr_selector2_134[15],addr_remain2_134[15:0],addr_remain2_134,addr_selector3_2159,addr_remain3_2159);


wire[15:0] addr_selector3_2160;
wire[15:0] addr_remain3_2160;
address_decode_4 decoder_3_2160 = address_decode_4(addr_selector2_135[0],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2160,addr_remain3_2160);


wire[15:0] addr_selector3_2161;
wire[15:0] addr_remain3_2161;
address_decode_4 decoder_3_2161 = address_decode_4(addr_selector2_135[1],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2161,addr_remain3_2161);


wire[15:0] addr_selector3_2162;
wire[15:0] addr_remain3_2162;
address_decode_4 decoder_3_2162 = address_decode_4(addr_selector2_135[2],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2162,addr_remain3_2162);


wire[15:0] addr_selector3_2163;
wire[15:0] addr_remain3_2163;
address_decode_4 decoder_3_2163 = address_decode_4(addr_selector2_135[3],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2163,addr_remain3_2163);


wire[15:0] addr_selector3_2164;
wire[15:0] addr_remain3_2164;
address_decode_4 decoder_3_2164 = address_decode_4(addr_selector2_135[4],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2164,addr_remain3_2164);


wire[15:0] addr_selector3_2165;
wire[15:0] addr_remain3_2165;
address_decode_4 decoder_3_2165 = address_decode_4(addr_selector2_135[5],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2165,addr_remain3_2165);


wire[15:0] addr_selector3_2166;
wire[15:0] addr_remain3_2166;
address_decode_4 decoder_3_2166 = address_decode_4(addr_selector2_135[6],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2166,addr_remain3_2166);


wire[15:0] addr_selector3_2167;
wire[15:0] addr_remain3_2167;
address_decode_4 decoder_3_2167 = address_decode_4(addr_selector2_135[7],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2167,addr_remain3_2167);


wire[15:0] addr_selector3_2168;
wire[15:0] addr_remain3_2168;
address_decode_4 decoder_3_2168 = address_decode_4(addr_selector2_135[8],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2168,addr_remain3_2168);


wire[15:0] addr_selector3_2169;
wire[15:0] addr_remain3_2169;
address_decode_4 decoder_3_2169 = address_decode_4(addr_selector2_135[9],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2169,addr_remain3_2169);


wire[15:0] addr_selector3_2170;
wire[15:0] addr_remain3_2170;
address_decode_4 decoder_3_2170 = address_decode_4(addr_selector2_135[10],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2170,addr_remain3_2170);


wire[15:0] addr_selector3_2171;
wire[15:0] addr_remain3_2171;
address_decode_4 decoder_3_2171 = address_decode_4(addr_selector2_135[11],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2171,addr_remain3_2171);


wire[15:0] addr_selector3_2172;
wire[15:0] addr_remain3_2172;
address_decode_4 decoder_3_2172 = address_decode_4(addr_selector2_135[12],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2172,addr_remain3_2172);


wire[15:0] addr_selector3_2173;
wire[15:0] addr_remain3_2173;
address_decode_4 decoder_3_2173 = address_decode_4(addr_selector2_135[13],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2173,addr_remain3_2173);


wire[15:0] addr_selector3_2174;
wire[15:0] addr_remain3_2174;
address_decode_4 decoder_3_2174 = address_decode_4(addr_selector2_135[14],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2174,addr_remain3_2174);


wire[15:0] addr_selector3_2175;
wire[15:0] addr_remain3_2175;
address_decode_4 decoder_3_2175 = address_decode_4(addr_selector2_135[15],addr_remain2_135[15:0],addr_remain2_135,addr_selector3_2175,addr_remain3_2175);


wire[15:0] addr_selector3_2176;
wire[15:0] addr_remain3_2176;
address_decode_4 decoder_3_2176 = address_decode_4(addr_selector2_136[0],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2176,addr_remain3_2176);


wire[15:0] addr_selector3_2177;
wire[15:0] addr_remain3_2177;
address_decode_4 decoder_3_2177 = address_decode_4(addr_selector2_136[1],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2177,addr_remain3_2177);


wire[15:0] addr_selector3_2178;
wire[15:0] addr_remain3_2178;
address_decode_4 decoder_3_2178 = address_decode_4(addr_selector2_136[2],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2178,addr_remain3_2178);


wire[15:0] addr_selector3_2179;
wire[15:0] addr_remain3_2179;
address_decode_4 decoder_3_2179 = address_decode_4(addr_selector2_136[3],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2179,addr_remain3_2179);


wire[15:0] addr_selector3_2180;
wire[15:0] addr_remain3_2180;
address_decode_4 decoder_3_2180 = address_decode_4(addr_selector2_136[4],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2180,addr_remain3_2180);


wire[15:0] addr_selector3_2181;
wire[15:0] addr_remain3_2181;
address_decode_4 decoder_3_2181 = address_decode_4(addr_selector2_136[5],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2181,addr_remain3_2181);


wire[15:0] addr_selector3_2182;
wire[15:0] addr_remain3_2182;
address_decode_4 decoder_3_2182 = address_decode_4(addr_selector2_136[6],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2182,addr_remain3_2182);


wire[15:0] addr_selector3_2183;
wire[15:0] addr_remain3_2183;
address_decode_4 decoder_3_2183 = address_decode_4(addr_selector2_136[7],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2183,addr_remain3_2183);


wire[15:0] addr_selector3_2184;
wire[15:0] addr_remain3_2184;
address_decode_4 decoder_3_2184 = address_decode_4(addr_selector2_136[8],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2184,addr_remain3_2184);


wire[15:0] addr_selector3_2185;
wire[15:0] addr_remain3_2185;
address_decode_4 decoder_3_2185 = address_decode_4(addr_selector2_136[9],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2185,addr_remain3_2185);


wire[15:0] addr_selector3_2186;
wire[15:0] addr_remain3_2186;
address_decode_4 decoder_3_2186 = address_decode_4(addr_selector2_136[10],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2186,addr_remain3_2186);


wire[15:0] addr_selector3_2187;
wire[15:0] addr_remain3_2187;
address_decode_4 decoder_3_2187 = address_decode_4(addr_selector2_136[11],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2187,addr_remain3_2187);


wire[15:0] addr_selector3_2188;
wire[15:0] addr_remain3_2188;
address_decode_4 decoder_3_2188 = address_decode_4(addr_selector2_136[12],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2188,addr_remain3_2188);


wire[15:0] addr_selector3_2189;
wire[15:0] addr_remain3_2189;
address_decode_4 decoder_3_2189 = address_decode_4(addr_selector2_136[13],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2189,addr_remain3_2189);


wire[15:0] addr_selector3_2190;
wire[15:0] addr_remain3_2190;
address_decode_4 decoder_3_2190 = address_decode_4(addr_selector2_136[14],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2190,addr_remain3_2190);


wire[15:0] addr_selector3_2191;
wire[15:0] addr_remain3_2191;
address_decode_4 decoder_3_2191 = address_decode_4(addr_selector2_136[15],addr_remain2_136[15:0],addr_remain2_136,addr_selector3_2191,addr_remain3_2191);


wire[15:0] addr_selector3_2192;
wire[15:0] addr_remain3_2192;
address_decode_4 decoder_3_2192 = address_decode_4(addr_selector2_137[0],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2192,addr_remain3_2192);


wire[15:0] addr_selector3_2193;
wire[15:0] addr_remain3_2193;
address_decode_4 decoder_3_2193 = address_decode_4(addr_selector2_137[1],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2193,addr_remain3_2193);


wire[15:0] addr_selector3_2194;
wire[15:0] addr_remain3_2194;
address_decode_4 decoder_3_2194 = address_decode_4(addr_selector2_137[2],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2194,addr_remain3_2194);


wire[15:0] addr_selector3_2195;
wire[15:0] addr_remain3_2195;
address_decode_4 decoder_3_2195 = address_decode_4(addr_selector2_137[3],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2195,addr_remain3_2195);


wire[15:0] addr_selector3_2196;
wire[15:0] addr_remain3_2196;
address_decode_4 decoder_3_2196 = address_decode_4(addr_selector2_137[4],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2196,addr_remain3_2196);


wire[15:0] addr_selector3_2197;
wire[15:0] addr_remain3_2197;
address_decode_4 decoder_3_2197 = address_decode_4(addr_selector2_137[5],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2197,addr_remain3_2197);


wire[15:0] addr_selector3_2198;
wire[15:0] addr_remain3_2198;
address_decode_4 decoder_3_2198 = address_decode_4(addr_selector2_137[6],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2198,addr_remain3_2198);


wire[15:0] addr_selector3_2199;
wire[15:0] addr_remain3_2199;
address_decode_4 decoder_3_2199 = address_decode_4(addr_selector2_137[7],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2199,addr_remain3_2199);


wire[15:0] addr_selector3_2200;
wire[15:0] addr_remain3_2200;
address_decode_4 decoder_3_2200 = address_decode_4(addr_selector2_137[8],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2200,addr_remain3_2200);


wire[15:0] addr_selector3_2201;
wire[15:0] addr_remain3_2201;
address_decode_4 decoder_3_2201 = address_decode_4(addr_selector2_137[9],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2201,addr_remain3_2201);


wire[15:0] addr_selector3_2202;
wire[15:0] addr_remain3_2202;
address_decode_4 decoder_3_2202 = address_decode_4(addr_selector2_137[10],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2202,addr_remain3_2202);


wire[15:0] addr_selector3_2203;
wire[15:0] addr_remain3_2203;
address_decode_4 decoder_3_2203 = address_decode_4(addr_selector2_137[11],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2203,addr_remain3_2203);


wire[15:0] addr_selector3_2204;
wire[15:0] addr_remain3_2204;
address_decode_4 decoder_3_2204 = address_decode_4(addr_selector2_137[12],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2204,addr_remain3_2204);


wire[15:0] addr_selector3_2205;
wire[15:0] addr_remain3_2205;
address_decode_4 decoder_3_2205 = address_decode_4(addr_selector2_137[13],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2205,addr_remain3_2205);


wire[15:0] addr_selector3_2206;
wire[15:0] addr_remain3_2206;
address_decode_4 decoder_3_2206 = address_decode_4(addr_selector2_137[14],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2206,addr_remain3_2206);


wire[15:0] addr_selector3_2207;
wire[15:0] addr_remain3_2207;
address_decode_4 decoder_3_2207 = address_decode_4(addr_selector2_137[15],addr_remain2_137[15:0],addr_remain2_137,addr_selector3_2207,addr_remain3_2207);


wire[15:0] addr_selector3_2208;
wire[15:0] addr_remain3_2208;
address_decode_4 decoder_3_2208 = address_decode_4(addr_selector2_138[0],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2208,addr_remain3_2208);


wire[15:0] addr_selector3_2209;
wire[15:0] addr_remain3_2209;
address_decode_4 decoder_3_2209 = address_decode_4(addr_selector2_138[1],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2209,addr_remain3_2209);


wire[15:0] addr_selector3_2210;
wire[15:0] addr_remain3_2210;
address_decode_4 decoder_3_2210 = address_decode_4(addr_selector2_138[2],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2210,addr_remain3_2210);


wire[15:0] addr_selector3_2211;
wire[15:0] addr_remain3_2211;
address_decode_4 decoder_3_2211 = address_decode_4(addr_selector2_138[3],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2211,addr_remain3_2211);


wire[15:0] addr_selector3_2212;
wire[15:0] addr_remain3_2212;
address_decode_4 decoder_3_2212 = address_decode_4(addr_selector2_138[4],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2212,addr_remain3_2212);


wire[15:0] addr_selector3_2213;
wire[15:0] addr_remain3_2213;
address_decode_4 decoder_3_2213 = address_decode_4(addr_selector2_138[5],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2213,addr_remain3_2213);


wire[15:0] addr_selector3_2214;
wire[15:0] addr_remain3_2214;
address_decode_4 decoder_3_2214 = address_decode_4(addr_selector2_138[6],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2214,addr_remain3_2214);


wire[15:0] addr_selector3_2215;
wire[15:0] addr_remain3_2215;
address_decode_4 decoder_3_2215 = address_decode_4(addr_selector2_138[7],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2215,addr_remain3_2215);


wire[15:0] addr_selector3_2216;
wire[15:0] addr_remain3_2216;
address_decode_4 decoder_3_2216 = address_decode_4(addr_selector2_138[8],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2216,addr_remain3_2216);


wire[15:0] addr_selector3_2217;
wire[15:0] addr_remain3_2217;
address_decode_4 decoder_3_2217 = address_decode_4(addr_selector2_138[9],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2217,addr_remain3_2217);


wire[15:0] addr_selector3_2218;
wire[15:0] addr_remain3_2218;
address_decode_4 decoder_3_2218 = address_decode_4(addr_selector2_138[10],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2218,addr_remain3_2218);


wire[15:0] addr_selector3_2219;
wire[15:0] addr_remain3_2219;
address_decode_4 decoder_3_2219 = address_decode_4(addr_selector2_138[11],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2219,addr_remain3_2219);


wire[15:0] addr_selector3_2220;
wire[15:0] addr_remain3_2220;
address_decode_4 decoder_3_2220 = address_decode_4(addr_selector2_138[12],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2220,addr_remain3_2220);


wire[15:0] addr_selector3_2221;
wire[15:0] addr_remain3_2221;
address_decode_4 decoder_3_2221 = address_decode_4(addr_selector2_138[13],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2221,addr_remain3_2221);


wire[15:0] addr_selector3_2222;
wire[15:0] addr_remain3_2222;
address_decode_4 decoder_3_2222 = address_decode_4(addr_selector2_138[14],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2222,addr_remain3_2222);


wire[15:0] addr_selector3_2223;
wire[15:0] addr_remain3_2223;
address_decode_4 decoder_3_2223 = address_decode_4(addr_selector2_138[15],addr_remain2_138[15:0],addr_remain2_138,addr_selector3_2223,addr_remain3_2223);


wire[15:0] addr_selector3_2224;
wire[15:0] addr_remain3_2224;
address_decode_4 decoder_3_2224 = address_decode_4(addr_selector2_139[0],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2224,addr_remain3_2224);


wire[15:0] addr_selector3_2225;
wire[15:0] addr_remain3_2225;
address_decode_4 decoder_3_2225 = address_decode_4(addr_selector2_139[1],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2225,addr_remain3_2225);


wire[15:0] addr_selector3_2226;
wire[15:0] addr_remain3_2226;
address_decode_4 decoder_3_2226 = address_decode_4(addr_selector2_139[2],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2226,addr_remain3_2226);


wire[15:0] addr_selector3_2227;
wire[15:0] addr_remain3_2227;
address_decode_4 decoder_3_2227 = address_decode_4(addr_selector2_139[3],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2227,addr_remain3_2227);


wire[15:0] addr_selector3_2228;
wire[15:0] addr_remain3_2228;
address_decode_4 decoder_3_2228 = address_decode_4(addr_selector2_139[4],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2228,addr_remain3_2228);


wire[15:0] addr_selector3_2229;
wire[15:0] addr_remain3_2229;
address_decode_4 decoder_3_2229 = address_decode_4(addr_selector2_139[5],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2229,addr_remain3_2229);


wire[15:0] addr_selector3_2230;
wire[15:0] addr_remain3_2230;
address_decode_4 decoder_3_2230 = address_decode_4(addr_selector2_139[6],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2230,addr_remain3_2230);


wire[15:0] addr_selector3_2231;
wire[15:0] addr_remain3_2231;
address_decode_4 decoder_3_2231 = address_decode_4(addr_selector2_139[7],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2231,addr_remain3_2231);


wire[15:0] addr_selector3_2232;
wire[15:0] addr_remain3_2232;
address_decode_4 decoder_3_2232 = address_decode_4(addr_selector2_139[8],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2232,addr_remain3_2232);


wire[15:0] addr_selector3_2233;
wire[15:0] addr_remain3_2233;
address_decode_4 decoder_3_2233 = address_decode_4(addr_selector2_139[9],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2233,addr_remain3_2233);


wire[15:0] addr_selector3_2234;
wire[15:0] addr_remain3_2234;
address_decode_4 decoder_3_2234 = address_decode_4(addr_selector2_139[10],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2234,addr_remain3_2234);


wire[15:0] addr_selector3_2235;
wire[15:0] addr_remain3_2235;
address_decode_4 decoder_3_2235 = address_decode_4(addr_selector2_139[11],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2235,addr_remain3_2235);


wire[15:0] addr_selector3_2236;
wire[15:0] addr_remain3_2236;
address_decode_4 decoder_3_2236 = address_decode_4(addr_selector2_139[12],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2236,addr_remain3_2236);


wire[15:0] addr_selector3_2237;
wire[15:0] addr_remain3_2237;
address_decode_4 decoder_3_2237 = address_decode_4(addr_selector2_139[13],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2237,addr_remain3_2237);


wire[15:0] addr_selector3_2238;
wire[15:0] addr_remain3_2238;
address_decode_4 decoder_3_2238 = address_decode_4(addr_selector2_139[14],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2238,addr_remain3_2238);


wire[15:0] addr_selector3_2239;
wire[15:0] addr_remain3_2239;
address_decode_4 decoder_3_2239 = address_decode_4(addr_selector2_139[15],addr_remain2_139[15:0],addr_remain2_139,addr_selector3_2239,addr_remain3_2239);


wire[15:0] addr_selector3_2240;
wire[15:0] addr_remain3_2240;
address_decode_4 decoder_3_2240 = address_decode_4(addr_selector2_140[0],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2240,addr_remain3_2240);


wire[15:0] addr_selector3_2241;
wire[15:0] addr_remain3_2241;
address_decode_4 decoder_3_2241 = address_decode_4(addr_selector2_140[1],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2241,addr_remain3_2241);


wire[15:0] addr_selector3_2242;
wire[15:0] addr_remain3_2242;
address_decode_4 decoder_3_2242 = address_decode_4(addr_selector2_140[2],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2242,addr_remain3_2242);


wire[15:0] addr_selector3_2243;
wire[15:0] addr_remain3_2243;
address_decode_4 decoder_3_2243 = address_decode_4(addr_selector2_140[3],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2243,addr_remain3_2243);


wire[15:0] addr_selector3_2244;
wire[15:0] addr_remain3_2244;
address_decode_4 decoder_3_2244 = address_decode_4(addr_selector2_140[4],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2244,addr_remain3_2244);


wire[15:0] addr_selector3_2245;
wire[15:0] addr_remain3_2245;
address_decode_4 decoder_3_2245 = address_decode_4(addr_selector2_140[5],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2245,addr_remain3_2245);


wire[15:0] addr_selector3_2246;
wire[15:0] addr_remain3_2246;
address_decode_4 decoder_3_2246 = address_decode_4(addr_selector2_140[6],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2246,addr_remain3_2246);


wire[15:0] addr_selector3_2247;
wire[15:0] addr_remain3_2247;
address_decode_4 decoder_3_2247 = address_decode_4(addr_selector2_140[7],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2247,addr_remain3_2247);


wire[15:0] addr_selector3_2248;
wire[15:0] addr_remain3_2248;
address_decode_4 decoder_3_2248 = address_decode_4(addr_selector2_140[8],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2248,addr_remain3_2248);


wire[15:0] addr_selector3_2249;
wire[15:0] addr_remain3_2249;
address_decode_4 decoder_3_2249 = address_decode_4(addr_selector2_140[9],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2249,addr_remain3_2249);


wire[15:0] addr_selector3_2250;
wire[15:0] addr_remain3_2250;
address_decode_4 decoder_3_2250 = address_decode_4(addr_selector2_140[10],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2250,addr_remain3_2250);


wire[15:0] addr_selector3_2251;
wire[15:0] addr_remain3_2251;
address_decode_4 decoder_3_2251 = address_decode_4(addr_selector2_140[11],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2251,addr_remain3_2251);


wire[15:0] addr_selector3_2252;
wire[15:0] addr_remain3_2252;
address_decode_4 decoder_3_2252 = address_decode_4(addr_selector2_140[12],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2252,addr_remain3_2252);


wire[15:0] addr_selector3_2253;
wire[15:0] addr_remain3_2253;
address_decode_4 decoder_3_2253 = address_decode_4(addr_selector2_140[13],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2253,addr_remain3_2253);


wire[15:0] addr_selector3_2254;
wire[15:0] addr_remain3_2254;
address_decode_4 decoder_3_2254 = address_decode_4(addr_selector2_140[14],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2254,addr_remain3_2254);


wire[15:0] addr_selector3_2255;
wire[15:0] addr_remain3_2255;
address_decode_4 decoder_3_2255 = address_decode_4(addr_selector2_140[15],addr_remain2_140[15:0],addr_remain2_140,addr_selector3_2255,addr_remain3_2255);


wire[15:0] addr_selector3_2256;
wire[15:0] addr_remain3_2256;
address_decode_4 decoder_3_2256 = address_decode_4(addr_selector2_141[0],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2256,addr_remain3_2256);


wire[15:0] addr_selector3_2257;
wire[15:0] addr_remain3_2257;
address_decode_4 decoder_3_2257 = address_decode_4(addr_selector2_141[1],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2257,addr_remain3_2257);


wire[15:0] addr_selector3_2258;
wire[15:0] addr_remain3_2258;
address_decode_4 decoder_3_2258 = address_decode_4(addr_selector2_141[2],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2258,addr_remain3_2258);


wire[15:0] addr_selector3_2259;
wire[15:0] addr_remain3_2259;
address_decode_4 decoder_3_2259 = address_decode_4(addr_selector2_141[3],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2259,addr_remain3_2259);


wire[15:0] addr_selector3_2260;
wire[15:0] addr_remain3_2260;
address_decode_4 decoder_3_2260 = address_decode_4(addr_selector2_141[4],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2260,addr_remain3_2260);


wire[15:0] addr_selector3_2261;
wire[15:0] addr_remain3_2261;
address_decode_4 decoder_3_2261 = address_decode_4(addr_selector2_141[5],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2261,addr_remain3_2261);


wire[15:0] addr_selector3_2262;
wire[15:0] addr_remain3_2262;
address_decode_4 decoder_3_2262 = address_decode_4(addr_selector2_141[6],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2262,addr_remain3_2262);


wire[15:0] addr_selector3_2263;
wire[15:0] addr_remain3_2263;
address_decode_4 decoder_3_2263 = address_decode_4(addr_selector2_141[7],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2263,addr_remain3_2263);


wire[15:0] addr_selector3_2264;
wire[15:0] addr_remain3_2264;
address_decode_4 decoder_3_2264 = address_decode_4(addr_selector2_141[8],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2264,addr_remain3_2264);


wire[15:0] addr_selector3_2265;
wire[15:0] addr_remain3_2265;
address_decode_4 decoder_3_2265 = address_decode_4(addr_selector2_141[9],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2265,addr_remain3_2265);


wire[15:0] addr_selector3_2266;
wire[15:0] addr_remain3_2266;
address_decode_4 decoder_3_2266 = address_decode_4(addr_selector2_141[10],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2266,addr_remain3_2266);


wire[15:0] addr_selector3_2267;
wire[15:0] addr_remain3_2267;
address_decode_4 decoder_3_2267 = address_decode_4(addr_selector2_141[11],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2267,addr_remain3_2267);


wire[15:0] addr_selector3_2268;
wire[15:0] addr_remain3_2268;
address_decode_4 decoder_3_2268 = address_decode_4(addr_selector2_141[12],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2268,addr_remain3_2268);


wire[15:0] addr_selector3_2269;
wire[15:0] addr_remain3_2269;
address_decode_4 decoder_3_2269 = address_decode_4(addr_selector2_141[13],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2269,addr_remain3_2269);


wire[15:0] addr_selector3_2270;
wire[15:0] addr_remain3_2270;
address_decode_4 decoder_3_2270 = address_decode_4(addr_selector2_141[14],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2270,addr_remain3_2270);


wire[15:0] addr_selector3_2271;
wire[15:0] addr_remain3_2271;
address_decode_4 decoder_3_2271 = address_decode_4(addr_selector2_141[15],addr_remain2_141[15:0],addr_remain2_141,addr_selector3_2271,addr_remain3_2271);


wire[15:0] addr_selector3_2272;
wire[15:0] addr_remain3_2272;
address_decode_4 decoder_3_2272 = address_decode_4(addr_selector2_142[0],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2272,addr_remain3_2272);


wire[15:0] addr_selector3_2273;
wire[15:0] addr_remain3_2273;
address_decode_4 decoder_3_2273 = address_decode_4(addr_selector2_142[1],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2273,addr_remain3_2273);


wire[15:0] addr_selector3_2274;
wire[15:0] addr_remain3_2274;
address_decode_4 decoder_3_2274 = address_decode_4(addr_selector2_142[2],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2274,addr_remain3_2274);


wire[15:0] addr_selector3_2275;
wire[15:0] addr_remain3_2275;
address_decode_4 decoder_3_2275 = address_decode_4(addr_selector2_142[3],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2275,addr_remain3_2275);


wire[15:0] addr_selector3_2276;
wire[15:0] addr_remain3_2276;
address_decode_4 decoder_3_2276 = address_decode_4(addr_selector2_142[4],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2276,addr_remain3_2276);


wire[15:0] addr_selector3_2277;
wire[15:0] addr_remain3_2277;
address_decode_4 decoder_3_2277 = address_decode_4(addr_selector2_142[5],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2277,addr_remain3_2277);


wire[15:0] addr_selector3_2278;
wire[15:0] addr_remain3_2278;
address_decode_4 decoder_3_2278 = address_decode_4(addr_selector2_142[6],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2278,addr_remain3_2278);


wire[15:0] addr_selector3_2279;
wire[15:0] addr_remain3_2279;
address_decode_4 decoder_3_2279 = address_decode_4(addr_selector2_142[7],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2279,addr_remain3_2279);


wire[15:0] addr_selector3_2280;
wire[15:0] addr_remain3_2280;
address_decode_4 decoder_3_2280 = address_decode_4(addr_selector2_142[8],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2280,addr_remain3_2280);


wire[15:0] addr_selector3_2281;
wire[15:0] addr_remain3_2281;
address_decode_4 decoder_3_2281 = address_decode_4(addr_selector2_142[9],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2281,addr_remain3_2281);


wire[15:0] addr_selector3_2282;
wire[15:0] addr_remain3_2282;
address_decode_4 decoder_3_2282 = address_decode_4(addr_selector2_142[10],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2282,addr_remain3_2282);


wire[15:0] addr_selector3_2283;
wire[15:0] addr_remain3_2283;
address_decode_4 decoder_3_2283 = address_decode_4(addr_selector2_142[11],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2283,addr_remain3_2283);


wire[15:0] addr_selector3_2284;
wire[15:0] addr_remain3_2284;
address_decode_4 decoder_3_2284 = address_decode_4(addr_selector2_142[12],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2284,addr_remain3_2284);


wire[15:0] addr_selector3_2285;
wire[15:0] addr_remain3_2285;
address_decode_4 decoder_3_2285 = address_decode_4(addr_selector2_142[13],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2285,addr_remain3_2285);


wire[15:0] addr_selector3_2286;
wire[15:0] addr_remain3_2286;
address_decode_4 decoder_3_2286 = address_decode_4(addr_selector2_142[14],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2286,addr_remain3_2286);


wire[15:0] addr_selector3_2287;
wire[15:0] addr_remain3_2287;
address_decode_4 decoder_3_2287 = address_decode_4(addr_selector2_142[15],addr_remain2_142[15:0],addr_remain2_142,addr_selector3_2287,addr_remain3_2287);


wire[15:0] addr_selector3_2288;
wire[15:0] addr_remain3_2288;
address_decode_4 decoder_3_2288 = address_decode_4(addr_selector2_143[0],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2288,addr_remain3_2288);


wire[15:0] addr_selector3_2289;
wire[15:0] addr_remain3_2289;
address_decode_4 decoder_3_2289 = address_decode_4(addr_selector2_143[1],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2289,addr_remain3_2289);


wire[15:0] addr_selector3_2290;
wire[15:0] addr_remain3_2290;
address_decode_4 decoder_3_2290 = address_decode_4(addr_selector2_143[2],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2290,addr_remain3_2290);


wire[15:0] addr_selector3_2291;
wire[15:0] addr_remain3_2291;
address_decode_4 decoder_3_2291 = address_decode_4(addr_selector2_143[3],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2291,addr_remain3_2291);


wire[15:0] addr_selector3_2292;
wire[15:0] addr_remain3_2292;
address_decode_4 decoder_3_2292 = address_decode_4(addr_selector2_143[4],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2292,addr_remain3_2292);


wire[15:0] addr_selector3_2293;
wire[15:0] addr_remain3_2293;
address_decode_4 decoder_3_2293 = address_decode_4(addr_selector2_143[5],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2293,addr_remain3_2293);


wire[15:0] addr_selector3_2294;
wire[15:0] addr_remain3_2294;
address_decode_4 decoder_3_2294 = address_decode_4(addr_selector2_143[6],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2294,addr_remain3_2294);


wire[15:0] addr_selector3_2295;
wire[15:0] addr_remain3_2295;
address_decode_4 decoder_3_2295 = address_decode_4(addr_selector2_143[7],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2295,addr_remain3_2295);


wire[15:0] addr_selector3_2296;
wire[15:0] addr_remain3_2296;
address_decode_4 decoder_3_2296 = address_decode_4(addr_selector2_143[8],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2296,addr_remain3_2296);


wire[15:0] addr_selector3_2297;
wire[15:0] addr_remain3_2297;
address_decode_4 decoder_3_2297 = address_decode_4(addr_selector2_143[9],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2297,addr_remain3_2297);


wire[15:0] addr_selector3_2298;
wire[15:0] addr_remain3_2298;
address_decode_4 decoder_3_2298 = address_decode_4(addr_selector2_143[10],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2298,addr_remain3_2298);


wire[15:0] addr_selector3_2299;
wire[15:0] addr_remain3_2299;
address_decode_4 decoder_3_2299 = address_decode_4(addr_selector2_143[11],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2299,addr_remain3_2299);


wire[15:0] addr_selector3_2300;
wire[15:0] addr_remain3_2300;
address_decode_4 decoder_3_2300 = address_decode_4(addr_selector2_143[12],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2300,addr_remain3_2300);


wire[15:0] addr_selector3_2301;
wire[15:0] addr_remain3_2301;
address_decode_4 decoder_3_2301 = address_decode_4(addr_selector2_143[13],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2301,addr_remain3_2301);


wire[15:0] addr_selector3_2302;
wire[15:0] addr_remain3_2302;
address_decode_4 decoder_3_2302 = address_decode_4(addr_selector2_143[14],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2302,addr_remain3_2302);


wire[15:0] addr_selector3_2303;
wire[15:0] addr_remain3_2303;
address_decode_4 decoder_3_2303 = address_decode_4(addr_selector2_143[15],addr_remain2_143[15:0],addr_remain2_143,addr_selector3_2303,addr_remain3_2303);


wire[15:0] addr_selector3_2304;
wire[15:0] addr_remain3_2304;
address_decode_4 decoder_3_2304 = address_decode_4(addr_selector2_144[0],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2304,addr_remain3_2304);


wire[15:0] addr_selector3_2305;
wire[15:0] addr_remain3_2305;
address_decode_4 decoder_3_2305 = address_decode_4(addr_selector2_144[1],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2305,addr_remain3_2305);


wire[15:0] addr_selector3_2306;
wire[15:0] addr_remain3_2306;
address_decode_4 decoder_3_2306 = address_decode_4(addr_selector2_144[2],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2306,addr_remain3_2306);


wire[15:0] addr_selector3_2307;
wire[15:0] addr_remain3_2307;
address_decode_4 decoder_3_2307 = address_decode_4(addr_selector2_144[3],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2307,addr_remain3_2307);


wire[15:0] addr_selector3_2308;
wire[15:0] addr_remain3_2308;
address_decode_4 decoder_3_2308 = address_decode_4(addr_selector2_144[4],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2308,addr_remain3_2308);


wire[15:0] addr_selector3_2309;
wire[15:0] addr_remain3_2309;
address_decode_4 decoder_3_2309 = address_decode_4(addr_selector2_144[5],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2309,addr_remain3_2309);


wire[15:0] addr_selector3_2310;
wire[15:0] addr_remain3_2310;
address_decode_4 decoder_3_2310 = address_decode_4(addr_selector2_144[6],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2310,addr_remain3_2310);


wire[15:0] addr_selector3_2311;
wire[15:0] addr_remain3_2311;
address_decode_4 decoder_3_2311 = address_decode_4(addr_selector2_144[7],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2311,addr_remain3_2311);


wire[15:0] addr_selector3_2312;
wire[15:0] addr_remain3_2312;
address_decode_4 decoder_3_2312 = address_decode_4(addr_selector2_144[8],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2312,addr_remain3_2312);


wire[15:0] addr_selector3_2313;
wire[15:0] addr_remain3_2313;
address_decode_4 decoder_3_2313 = address_decode_4(addr_selector2_144[9],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2313,addr_remain3_2313);


wire[15:0] addr_selector3_2314;
wire[15:0] addr_remain3_2314;
address_decode_4 decoder_3_2314 = address_decode_4(addr_selector2_144[10],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2314,addr_remain3_2314);


wire[15:0] addr_selector3_2315;
wire[15:0] addr_remain3_2315;
address_decode_4 decoder_3_2315 = address_decode_4(addr_selector2_144[11],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2315,addr_remain3_2315);


wire[15:0] addr_selector3_2316;
wire[15:0] addr_remain3_2316;
address_decode_4 decoder_3_2316 = address_decode_4(addr_selector2_144[12],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2316,addr_remain3_2316);


wire[15:0] addr_selector3_2317;
wire[15:0] addr_remain3_2317;
address_decode_4 decoder_3_2317 = address_decode_4(addr_selector2_144[13],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2317,addr_remain3_2317);


wire[15:0] addr_selector3_2318;
wire[15:0] addr_remain3_2318;
address_decode_4 decoder_3_2318 = address_decode_4(addr_selector2_144[14],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2318,addr_remain3_2318);


wire[15:0] addr_selector3_2319;
wire[15:0] addr_remain3_2319;
address_decode_4 decoder_3_2319 = address_decode_4(addr_selector2_144[15],addr_remain2_144[15:0],addr_remain2_144,addr_selector3_2319,addr_remain3_2319);


wire[15:0] addr_selector3_2320;
wire[15:0] addr_remain3_2320;
address_decode_4 decoder_3_2320 = address_decode_4(addr_selector2_145[0],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2320,addr_remain3_2320);


wire[15:0] addr_selector3_2321;
wire[15:0] addr_remain3_2321;
address_decode_4 decoder_3_2321 = address_decode_4(addr_selector2_145[1],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2321,addr_remain3_2321);


wire[15:0] addr_selector3_2322;
wire[15:0] addr_remain3_2322;
address_decode_4 decoder_3_2322 = address_decode_4(addr_selector2_145[2],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2322,addr_remain3_2322);


wire[15:0] addr_selector3_2323;
wire[15:0] addr_remain3_2323;
address_decode_4 decoder_3_2323 = address_decode_4(addr_selector2_145[3],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2323,addr_remain3_2323);


wire[15:0] addr_selector3_2324;
wire[15:0] addr_remain3_2324;
address_decode_4 decoder_3_2324 = address_decode_4(addr_selector2_145[4],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2324,addr_remain3_2324);


wire[15:0] addr_selector3_2325;
wire[15:0] addr_remain3_2325;
address_decode_4 decoder_3_2325 = address_decode_4(addr_selector2_145[5],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2325,addr_remain3_2325);


wire[15:0] addr_selector3_2326;
wire[15:0] addr_remain3_2326;
address_decode_4 decoder_3_2326 = address_decode_4(addr_selector2_145[6],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2326,addr_remain3_2326);


wire[15:0] addr_selector3_2327;
wire[15:0] addr_remain3_2327;
address_decode_4 decoder_3_2327 = address_decode_4(addr_selector2_145[7],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2327,addr_remain3_2327);


wire[15:0] addr_selector3_2328;
wire[15:0] addr_remain3_2328;
address_decode_4 decoder_3_2328 = address_decode_4(addr_selector2_145[8],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2328,addr_remain3_2328);


wire[15:0] addr_selector3_2329;
wire[15:0] addr_remain3_2329;
address_decode_4 decoder_3_2329 = address_decode_4(addr_selector2_145[9],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2329,addr_remain3_2329);


wire[15:0] addr_selector3_2330;
wire[15:0] addr_remain3_2330;
address_decode_4 decoder_3_2330 = address_decode_4(addr_selector2_145[10],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2330,addr_remain3_2330);


wire[15:0] addr_selector3_2331;
wire[15:0] addr_remain3_2331;
address_decode_4 decoder_3_2331 = address_decode_4(addr_selector2_145[11],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2331,addr_remain3_2331);


wire[15:0] addr_selector3_2332;
wire[15:0] addr_remain3_2332;
address_decode_4 decoder_3_2332 = address_decode_4(addr_selector2_145[12],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2332,addr_remain3_2332);


wire[15:0] addr_selector3_2333;
wire[15:0] addr_remain3_2333;
address_decode_4 decoder_3_2333 = address_decode_4(addr_selector2_145[13],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2333,addr_remain3_2333);


wire[15:0] addr_selector3_2334;
wire[15:0] addr_remain3_2334;
address_decode_4 decoder_3_2334 = address_decode_4(addr_selector2_145[14],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2334,addr_remain3_2334);


wire[15:0] addr_selector3_2335;
wire[15:0] addr_remain3_2335;
address_decode_4 decoder_3_2335 = address_decode_4(addr_selector2_145[15],addr_remain2_145[15:0],addr_remain2_145,addr_selector3_2335,addr_remain3_2335);


wire[15:0] addr_selector3_2336;
wire[15:0] addr_remain3_2336;
address_decode_4 decoder_3_2336 = address_decode_4(addr_selector2_146[0],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2336,addr_remain3_2336);


wire[15:0] addr_selector3_2337;
wire[15:0] addr_remain3_2337;
address_decode_4 decoder_3_2337 = address_decode_4(addr_selector2_146[1],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2337,addr_remain3_2337);


wire[15:0] addr_selector3_2338;
wire[15:0] addr_remain3_2338;
address_decode_4 decoder_3_2338 = address_decode_4(addr_selector2_146[2],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2338,addr_remain3_2338);


wire[15:0] addr_selector3_2339;
wire[15:0] addr_remain3_2339;
address_decode_4 decoder_3_2339 = address_decode_4(addr_selector2_146[3],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2339,addr_remain3_2339);


wire[15:0] addr_selector3_2340;
wire[15:0] addr_remain3_2340;
address_decode_4 decoder_3_2340 = address_decode_4(addr_selector2_146[4],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2340,addr_remain3_2340);


wire[15:0] addr_selector3_2341;
wire[15:0] addr_remain3_2341;
address_decode_4 decoder_3_2341 = address_decode_4(addr_selector2_146[5],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2341,addr_remain3_2341);


wire[15:0] addr_selector3_2342;
wire[15:0] addr_remain3_2342;
address_decode_4 decoder_3_2342 = address_decode_4(addr_selector2_146[6],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2342,addr_remain3_2342);


wire[15:0] addr_selector3_2343;
wire[15:0] addr_remain3_2343;
address_decode_4 decoder_3_2343 = address_decode_4(addr_selector2_146[7],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2343,addr_remain3_2343);


wire[15:0] addr_selector3_2344;
wire[15:0] addr_remain3_2344;
address_decode_4 decoder_3_2344 = address_decode_4(addr_selector2_146[8],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2344,addr_remain3_2344);


wire[15:0] addr_selector3_2345;
wire[15:0] addr_remain3_2345;
address_decode_4 decoder_3_2345 = address_decode_4(addr_selector2_146[9],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2345,addr_remain3_2345);


wire[15:0] addr_selector3_2346;
wire[15:0] addr_remain3_2346;
address_decode_4 decoder_3_2346 = address_decode_4(addr_selector2_146[10],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2346,addr_remain3_2346);


wire[15:0] addr_selector3_2347;
wire[15:0] addr_remain3_2347;
address_decode_4 decoder_3_2347 = address_decode_4(addr_selector2_146[11],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2347,addr_remain3_2347);


wire[15:0] addr_selector3_2348;
wire[15:0] addr_remain3_2348;
address_decode_4 decoder_3_2348 = address_decode_4(addr_selector2_146[12],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2348,addr_remain3_2348);


wire[15:0] addr_selector3_2349;
wire[15:0] addr_remain3_2349;
address_decode_4 decoder_3_2349 = address_decode_4(addr_selector2_146[13],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2349,addr_remain3_2349);


wire[15:0] addr_selector3_2350;
wire[15:0] addr_remain3_2350;
address_decode_4 decoder_3_2350 = address_decode_4(addr_selector2_146[14],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2350,addr_remain3_2350);


wire[15:0] addr_selector3_2351;
wire[15:0] addr_remain3_2351;
address_decode_4 decoder_3_2351 = address_decode_4(addr_selector2_146[15],addr_remain2_146[15:0],addr_remain2_146,addr_selector3_2351,addr_remain3_2351);


wire[15:0] addr_selector3_2352;
wire[15:0] addr_remain3_2352;
address_decode_4 decoder_3_2352 = address_decode_4(addr_selector2_147[0],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2352,addr_remain3_2352);


wire[15:0] addr_selector3_2353;
wire[15:0] addr_remain3_2353;
address_decode_4 decoder_3_2353 = address_decode_4(addr_selector2_147[1],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2353,addr_remain3_2353);


wire[15:0] addr_selector3_2354;
wire[15:0] addr_remain3_2354;
address_decode_4 decoder_3_2354 = address_decode_4(addr_selector2_147[2],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2354,addr_remain3_2354);


wire[15:0] addr_selector3_2355;
wire[15:0] addr_remain3_2355;
address_decode_4 decoder_3_2355 = address_decode_4(addr_selector2_147[3],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2355,addr_remain3_2355);


wire[15:0] addr_selector3_2356;
wire[15:0] addr_remain3_2356;
address_decode_4 decoder_3_2356 = address_decode_4(addr_selector2_147[4],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2356,addr_remain3_2356);


wire[15:0] addr_selector3_2357;
wire[15:0] addr_remain3_2357;
address_decode_4 decoder_3_2357 = address_decode_4(addr_selector2_147[5],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2357,addr_remain3_2357);


wire[15:0] addr_selector3_2358;
wire[15:0] addr_remain3_2358;
address_decode_4 decoder_3_2358 = address_decode_4(addr_selector2_147[6],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2358,addr_remain3_2358);


wire[15:0] addr_selector3_2359;
wire[15:0] addr_remain3_2359;
address_decode_4 decoder_3_2359 = address_decode_4(addr_selector2_147[7],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2359,addr_remain3_2359);


wire[15:0] addr_selector3_2360;
wire[15:0] addr_remain3_2360;
address_decode_4 decoder_3_2360 = address_decode_4(addr_selector2_147[8],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2360,addr_remain3_2360);


wire[15:0] addr_selector3_2361;
wire[15:0] addr_remain3_2361;
address_decode_4 decoder_3_2361 = address_decode_4(addr_selector2_147[9],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2361,addr_remain3_2361);


wire[15:0] addr_selector3_2362;
wire[15:0] addr_remain3_2362;
address_decode_4 decoder_3_2362 = address_decode_4(addr_selector2_147[10],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2362,addr_remain3_2362);


wire[15:0] addr_selector3_2363;
wire[15:0] addr_remain3_2363;
address_decode_4 decoder_3_2363 = address_decode_4(addr_selector2_147[11],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2363,addr_remain3_2363);


wire[15:0] addr_selector3_2364;
wire[15:0] addr_remain3_2364;
address_decode_4 decoder_3_2364 = address_decode_4(addr_selector2_147[12],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2364,addr_remain3_2364);


wire[15:0] addr_selector3_2365;
wire[15:0] addr_remain3_2365;
address_decode_4 decoder_3_2365 = address_decode_4(addr_selector2_147[13],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2365,addr_remain3_2365);


wire[15:0] addr_selector3_2366;
wire[15:0] addr_remain3_2366;
address_decode_4 decoder_3_2366 = address_decode_4(addr_selector2_147[14],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2366,addr_remain3_2366);


wire[15:0] addr_selector3_2367;
wire[15:0] addr_remain3_2367;
address_decode_4 decoder_3_2367 = address_decode_4(addr_selector2_147[15],addr_remain2_147[15:0],addr_remain2_147,addr_selector3_2367,addr_remain3_2367);


wire[15:0] addr_selector3_2368;
wire[15:0] addr_remain3_2368;
address_decode_4 decoder_3_2368 = address_decode_4(addr_selector2_148[0],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2368,addr_remain3_2368);


wire[15:0] addr_selector3_2369;
wire[15:0] addr_remain3_2369;
address_decode_4 decoder_3_2369 = address_decode_4(addr_selector2_148[1],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2369,addr_remain3_2369);


wire[15:0] addr_selector3_2370;
wire[15:0] addr_remain3_2370;
address_decode_4 decoder_3_2370 = address_decode_4(addr_selector2_148[2],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2370,addr_remain3_2370);


wire[15:0] addr_selector3_2371;
wire[15:0] addr_remain3_2371;
address_decode_4 decoder_3_2371 = address_decode_4(addr_selector2_148[3],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2371,addr_remain3_2371);


wire[15:0] addr_selector3_2372;
wire[15:0] addr_remain3_2372;
address_decode_4 decoder_3_2372 = address_decode_4(addr_selector2_148[4],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2372,addr_remain3_2372);


wire[15:0] addr_selector3_2373;
wire[15:0] addr_remain3_2373;
address_decode_4 decoder_3_2373 = address_decode_4(addr_selector2_148[5],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2373,addr_remain3_2373);


wire[15:0] addr_selector3_2374;
wire[15:0] addr_remain3_2374;
address_decode_4 decoder_3_2374 = address_decode_4(addr_selector2_148[6],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2374,addr_remain3_2374);


wire[15:0] addr_selector3_2375;
wire[15:0] addr_remain3_2375;
address_decode_4 decoder_3_2375 = address_decode_4(addr_selector2_148[7],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2375,addr_remain3_2375);


wire[15:0] addr_selector3_2376;
wire[15:0] addr_remain3_2376;
address_decode_4 decoder_3_2376 = address_decode_4(addr_selector2_148[8],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2376,addr_remain3_2376);


wire[15:0] addr_selector3_2377;
wire[15:0] addr_remain3_2377;
address_decode_4 decoder_3_2377 = address_decode_4(addr_selector2_148[9],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2377,addr_remain3_2377);


wire[15:0] addr_selector3_2378;
wire[15:0] addr_remain3_2378;
address_decode_4 decoder_3_2378 = address_decode_4(addr_selector2_148[10],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2378,addr_remain3_2378);


wire[15:0] addr_selector3_2379;
wire[15:0] addr_remain3_2379;
address_decode_4 decoder_3_2379 = address_decode_4(addr_selector2_148[11],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2379,addr_remain3_2379);


wire[15:0] addr_selector3_2380;
wire[15:0] addr_remain3_2380;
address_decode_4 decoder_3_2380 = address_decode_4(addr_selector2_148[12],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2380,addr_remain3_2380);


wire[15:0] addr_selector3_2381;
wire[15:0] addr_remain3_2381;
address_decode_4 decoder_3_2381 = address_decode_4(addr_selector2_148[13],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2381,addr_remain3_2381);


wire[15:0] addr_selector3_2382;
wire[15:0] addr_remain3_2382;
address_decode_4 decoder_3_2382 = address_decode_4(addr_selector2_148[14],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2382,addr_remain3_2382);


wire[15:0] addr_selector3_2383;
wire[15:0] addr_remain3_2383;
address_decode_4 decoder_3_2383 = address_decode_4(addr_selector2_148[15],addr_remain2_148[15:0],addr_remain2_148,addr_selector3_2383,addr_remain3_2383);


wire[15:0] addr_selector3_2384;
wire[15:0] addr_remain3_2384;
address_decode_4 decoder_3_2384 = address_decode_4(addr_selector2_149[0],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2384,addr_remain3_2384);


wire[15:0] addr_selector3_2385;
wire[15:0] addr_remain3_2385;
address_decode_4 decoder_3_2385 = address_decode_4(addr_selector2_149[1],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2385,addr_remain3_2385);


wire[15:0] addr_selector3_2386;
wire[15:0] addr_remain3_2386;
address_decode_4 decoder_3_2386 = address_decode_4(addr_selector2_149[2],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2386,addr_remain3_2386);


wire[15:0] addr_selector3_2387;
wire[15:0] addr_remain3_2387;
address_decode_4 decoder_3_2387 = address_decode_4(addr_selector2_149[3],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2387,addr_remain3_2387);


wire[15:0] addr_selector3_2388;
wire[15:0] addr_remain3_2388;
address_decode_4 decoder_3_2388 = address_decode_4(addr_selector2_149[4],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2388,addr_remain3_2388);


wire[15:0] addr_selector3_2389;
wire[15:0] addr_remain3_2389;
address_decode_4 decoder_3_2389 = address_decode_4(addr_selector2_149[5],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2389,addr_remain3_2389);


wire[15:0] addr_selector3_2390;
wire[15:0] addr_remain3_2390;
address_decode_4 decoder_3_2390 = address_decode_4(addr_selector2_149[6],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2390,addr_remain3_2390);


wire[15:0] addr_selector3_2391;
wire[15:0] addr_remain3_2391;
address_decode_4 decoder_3_2391 = address_decode_4(addr_selector2_149[7],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2391,addr_remain3_2391);


wire[15:0] addr_selector3_2392;
wire[15:0] addr_remain3_2392;
address_decode_4 decoder_3_2392 = address_decode_4(addr_selector2_149[8],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2392,addr_remain3_2392);


wire[15:0] addr_selector3_2393;
wire[15:0] addr_remain3_2393;
address_decode_4 decoder_3_2393 = address_decode_4(addr_selector2_149[9],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2393,addr_remain3_2393);


wire[15:0] addr_selector3_2394;
wire[15:0] addr_remain3_2394;
address_decode_4 decoder_3_2394 = address_decode_4(addr_selector2_149[10],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2394,addr_remain3_2394);


wire[15:0] addr_selector3_2395;
wire[15:0] addr_remain3_2395;
address_decode_4 decoder_3_2395 = address_decode_4(addr_selector2_149[11],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2395,addr_remain3_2395);


wire[15:0] addr_selector3_2396;
wire[15:0] addr_remain3_2396;
address_decode_4 decoder_3_2396 = address_decode_4(addr_selector2_149[12],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2396,addr_remain3_2396);


wire[15:0] addr_selector3_2397;
wire[15:0] addr_remain3_2397;
address_decode_4 decoder_3_2397 = address_decode_4(addr_selector2_149[13],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2397,addr_remain3_2397);


wire[15:0] addr_selector3_2398;
wire[15:0] addr_remain3_2398;
address_decode_4 decoder_3_2398 = address_decode_4(addr_selector2_149[14],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2398,addr_remain3_2398);


wire[15:0] addr_selector3_2399;
wire[15:0] addr_remain3_2399;
address_decode_4 decoder_3_2399 = address_decode_4(addr_selector2_149[15],addr_remain2_149[15:0],addr_remain2_149,addr_selector3_2399,addr_remain3_2399);


wire[15:0] addr_selector3_2400;
wire[15:0] addr_remain3_2400;
address_decode_4 decoder_3_2400 = address_decode_4(addr_selector2_150[0],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2400,addr_remain3_2400);


wire[15:0] addr_selector3_2401;
wire[15:0] addr_remain3_2401;
address_decode_4 decoder_3_2401 = address_decode_4(addr_selector2_150[1],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2401,addr_remain3_2401);


wire[15:0] addr_selector3_2402;
wire[15:0] addr_remain3_2402;
address_decode_4 decoder_3_2402 = address_decode_4(addr_selector2_150[2],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2402,addr_remain3_2402);


wire[15:0] addr_selector3_2403;
wire[15:0] addr_remain3_2403;
address_decode_4 decoder_3_2403 = address_decode_4(addr_selector2_150[3],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2403,addr_remain3_2403);


wire[15:0] addr_selector3_2404;
wire[15:0] addr_remain3_2404;
address_decode_4 decoder_3_2404 = address_decode_4(addr_selector2_150[4],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2404,addr_remain3_2404);


wire[15:0] addr_selector3_2405;
wire[15:0] addr_remain3_2405;
address_decode_4 decoder_3_2405 = address_decode_4(addr_selector2_150[5],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2405,addr_remain3_2405);


wire[15:0] addr_selector3_2406;
wire[15:0] addr_remain3_2406;
address_decode_4 decoder_3_2406 = address_decode_4(addr_selector2_150[6],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2406,addr_remain3_2406);


wire[15:0] addr_selector3_2407;
wire[15:0] addr_remain3_2407;
address_decode_4 decoder_3_2407 = address_decode_4(addr_selector2_150[7],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2407,addr_remain3_2407);


wire[15:0] addr_selector3_2408;
wire[15:0] addr_remain3_2408;
address_decode_4 decoder_3_2408 = address_decode_4(addr_selector2_150[8],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2408,addr_remain3_2408);


wire[15:0] addr_selector3_2409;
wire[15:0] addr_remain3_2409;
address_decode_4 decoder_3_2409 = address_decode_4(addr_selector2_150[9],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2409,addr_remain3_2409);


wire[15:0] addr_selector3_2410;
wire[15:0] addr_remain3_2410;
address_decode_4 decoder_3_2410 = address_decode_4(addr_selector2_150[10],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2410,addr_remain3_2410);


wire[15:0] addr_selector3_2411;
wire[15:0] addr_remain3_2411;
address_decode_4 decoder_3_2411 = address_decode_4(addr_selector2_150[11],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2411,addr_remain3_2411);


wire[15:0] addr_selector3_2412;
wire[15:0] addr_remain3_2412;
address_decode_4 decoder_3_2412 = address_decode_4(addr_selector2_150[12],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2412,addr_remain3_2412);


wire[15:0] addr_selector3_2413;
wire[15:0] addr_remain3_2413;
address_decode_4 decoder_3_2413 = address_decode_4(addr_selector2_150[13],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2413,addr_remain3_2413);


wire[15:0] addr_selector3_2414;
wire[15:0] addr_remain3_2414;
address_decode_4 decoder_3_2414 = address_decode_4(addr_selector2_150[14],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2414,addr_remain3_2414);


wire[15:0] addr_selector3_2415;
wire[15:0] addr_remain3_2415;
address_decode_4 decoder_3_2415 = address_decode_4(addr_selector2_150[15],addr_remain2_150[15:0],addr_remain2_150,addr_selector3_2415,addr_remain3_2415);


wire[15:0] addr_selector3_2416;
wire[15:0] addr_remain3_2416;
address_decode_4 decoder_3_2416 = address_decode_4(addr_selector2_151[0],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2416,addr_remain3_2416);


wire[15:0] addr_selector3_2417;
wire[15:0] addr_remain3_2417;
address_decode_4 decoder_3_2417 = address_decode_4(addr_selector2_151[1],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2417,addr_remain3_2417);


wire[15:0] addr_selector3_2418;
wire[15:0] addr_remain3_2418;
address_decode_4 decoder_3_2418 = address_decode_4(addr_selector2_151[2],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2418,addr_remain3_2418);


wire[15:0] addr_selector3_2419;
wire[15:0] addr_remain3_2419;
address_decode_4 decoder_3_2419 = address_decode_4(addr_selector2_151[3],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2419,addr_remain3_2419);


wire[15:0] addr_selector3_2420;
wire[15:0] addr_remain3_2420;
address_decode_4 decoder_3_2420 = address_decode_4(addr_selector2_151[4],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2420,addr_remain3_2420);


wire[15:0] addr_selector3_2421;
wire[15:0] addr_remain3_2421;
address_decode_4 decoder_3_2421 = address_decode_4(addr_selector2_151[5],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2421,addr_remain3_2421);


wire[15:0] addr_selector3_2422;
wire[15:0] addr_remain3_2422;
address_decode_4 decoder_3_2422 = address_decode_4(addr_selector2_151[6],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2422,addr_remain3_2422);


wire[15:0] addr_selector3_2423;
wire[15:0] addr_remain3_2423;
address_decode_4 decoder_3_2423 = address_decode_4(addr_selector2_151[7],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2423,addr_remain3_2423);


wire[15:0] addr_selector3_2424;
wire[15:0] addr_remain3_2424;
address_decode_4 decoder_3_2424 = address_decode_4(addr_selector2_151[8],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2424,addr_remain3_2424);


wire[15:0] addr_selector3_2425;
wire[15:0] addr_remain3_2425;
address_decode_4 decoder_3_2425 = address_decode_4(addr_selector2_151[9],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2425,addr_remain3_2425);


wire[15:0] addr_selector3_2426;
wire[15:0] addr_remain3_2426;
address_decode_4 decoder_3_2426 = address_decode_4(addr_selector2_151[10],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2426,addr_remain3_2426);


wire[15:0] addr_selector3_2427;
wire[15:0] addr_remain3_2427;
address_decode_4 decoder_3_2427 = address_decode_4(addr_selector2_151[11],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2427,addr_remain3_2427);


wire[15:0] addr_selector3_2428;
wire[15:0] addr_remain3_2428;
address_decode_4 decoder_3_2428 = address_decode_4(addr_selector2_151[12],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2428,addr_remain3_2428);


wire[15:0] addr_selector3_2429;
wire[15:0] addr_remain3_2429;
address_decode_4 decoder_3_2429 = address_decode_4(addr_selector2_151[13],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2429,addr_remain3_2429);


wire[15:0] addr_selector3_2430;
wire[15:0] addr_remain3_2430;
address_decode_4 decoder_3_2430 = address_decode_4(addr_selector2_151[14],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2430,addr_remain3_2430);


wire[15:0] addr_selector3_2431;
wire[15:0] addr_remain3_2431;
address_decode_4 decoder_3_2431 = address_decode_4(addr_selector2_151[15],addr_remain2_151[15:0],addr_remain2_151,addr_selector3_2431,addr_remain3_2431);


wire[15:0] addr_selector3_2432;
wire[15:0] addr_remain3_2432;
address_decode_4 decoder_3_2432 = address_decode_4(addr_selector2_152[0],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2432,addr_remain3_2432);


wire[15:0] addr_selector3_2433;
wire[15:0] addr_remain3_2433;
address_decode_4 decoder_3_2433 = address_decode_4(addr_selector2_152[1],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2433,addr_remain3_2433);


wire[15:0] addr_selector3_2434;
wire[15:0] addr_remain3_2434;
address_decode_4 decoder_3_2434 = address_decode_4(addr_selector2_152[2],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2434,addr_remain3_2434);


wire[15:0] addr_selector3_2435;
wire[15:0] addr_remain3_2435;
address_decode_4 decoder_3_2435 = address_decode_4(addr_selector2_152[3],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2435,addr_remain3_2435);


wire[15:0] addr_selector3_2436;
wire[15:0] addr_remain3_2436;
address_decode_4 decoder_3_2436 = address_decode_4(addr_selector2_152[4],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2436,addr_remain3_2436);


wire[15:0] addr_selector3_2437;
wire[15:0] addr_remain3_2437;
address_decode_4 decoder_3_2437 = address_decode_4(addr_selector2_152[5],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2437,addr_remain3_2437);


wire[15:0] addr_selector3_2438;
wire[15:0] addr_remain3_2438;
address_decode_4 decoder_3_2438 = address_decode_4(addr_selector2_152[6],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2438,addr_remain3_2438);


wire[15:0] addr_selector3_2439;
wire[15:0] addr_remain3_2439;
address_decode_4 decoder_3_2439 = address_decode_4(addr_selector2_152[7],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2439,addr_remain3_2439);


wire[15:0] addr_selector3_2440;
wire[15:0] addr_remain3_2440;
address_decode_4 decoder_3_2440 = address_decode_4(addr_selector2_152[8],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2440,addr_remain3_2440);


wire[15:0] addr_selector3_2441;
wire[15:0] addr_remain3_2441;
address_decode_4 decoder_3_2441 = address_decode_4(addr_selector2_152[9],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2441,addr_remain3_2441);


wire[15:0] addr_selector3_2442;
wire[15:0] addr_remain3_2442;
address_decode_4 decoder_3_2442 = address_decode_4(addr_selector2_152[10],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2442,addr_remain3_2442);


wire[15:0] addr_selector3_2443;
wire[15:0] addr_remain3_2443;
address_decode_4 decoder_3_2443 = address_decode_4(addr_selector2_152[11],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2443,addr_remain3_2443);


wire[15:0] addr_selector3_2444;
wire[15:0] addr_remain3_2444;
address_decode_4 decoder_3_2444 = address_decode_4(addr_selector2_152[12],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2444,addr_remain3_2444);


wire[15:0] addr_selector3_2445;
wire[15:0] addr_remain3_2445;
address_decode_4 decoder_3_2445 = address_decode_4(addr_selector2_152[13],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2445,addr_remain3_2445);


wire[15:0] addr_selector3_2446;
wire[15:0] addr_remain3_2446;
address_decode_4 decoder_3_2446 = address_decode_4(addr_selector2_152[14],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2446,addr_remain3_2446);


wire[15:0] addr_selector3_2447;
wire[15:0] addr_remain3_2447;
address_decode_4 decoder_3_2447 = address_decode_4(addr_selector2_152[15],addr_remain2_152[15:0],addr_remain2_152,addr_selector3_2447,addr_remain3_2447);


wire[15:0] addr_selector3_2448;
wire[15:0] addr_remain3_2448;
address_decode_4 decoder_3_2448 = address_decode_4(addr_selector2_153[0],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2448,addr_remain3_2448);


wire[15:0] addr_selector3_2449;
wire[15:0] addr_remain3_2449;
address_decode_4 decoder_3_2449 = address_decode_4(addr_selector2_153[1],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2449,addr_remain3_2449);


wire[15:0] addr_selector3_2450;
wire[15:0] addr_remain3_2450;
address_decode_4 decoder_3_2450 = address_decode_4(addr_selector2_153[2],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2450,addr_remain3_2450);


wire[15:0] addr_selector3_2451;
wire[15:0] addr_remain3_2451;
address_decode_4 decoder_3_2451 = address_decode_4(addr_selector2_153[3],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2451,addr_remain3_2451);


wire[15:0] addr_selector3_2452;
wire[15:0] addr_remain3_2452;
address_decode_4 decoder_3_2452 = address_decode_4(addr_selector2_153[4],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2452,addr_remain3_2452);


wire[15:0] addr_selector3_2453;
wire[15:0] addr_remain3_2453;
address_decode_4 decoder_3_2453 = address_decode_4(addr_selector2_153[5],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2453,addr_remain3_2453);


wire[15:0] addr_selector3_2454;
wire[15:0] addr_remain3_2454;
address_decode_4 decoder_3_2454 = address_decode_4(addr_selector2_153[6],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2454,addr_remain3_2454);


wire[15:0] addr_selector3_2455;
wire[15:0] addr_remain3_2455;
address_decode_4 decoder_3_2455 = address_decode_4(addr_selector2_153[7],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2455,addr_remain3_2455);


wire[15:0] addr_selector3_2456;
wire[15:0] addr_remain3_2456;
address_decode_4 decoder_3_2456 = address_decode_4(addr_selector2_153[8],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2456,addr_remain3_2456);


wire[15:0] addr_selector3_2457;
wire[15:0] addr_remain3_2457;
address_decode_4 decoder_3_2457 = address_decode_4(addr_selector2_153[9],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2457,addr_remain3_2457);


wire[15:0] addr_selector3_2458;
wire[15:0] addr_remain3_2458;
address_decode_4 decoder_3_2458 = address_decode_4(addr_selector2_153[10],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2458,addr_remain3_2458);


wire[15:0] addr_selector3_2459;
wire[15:0] addr_remain3_2459;
address_decode_4 decoder_3_2459 = address_decode_4(addr_selector2_153[11],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2459,addr_remain3_2459);


wire[15:0] addr_selector3_2460;
wire[15:0] addr_remain3_2460;
address_decode_4 decoder_3_2460 = address_decode_4(addr_selector2_153[12],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2460,addr_remain3_2460);


wire[15:0] addr_selector3_2461;
wire[15:0] addr_remain3_2461;
address_decode_4 decoder_3_2461 = address_decode_4(addr_selector2_153[13],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2461,addr_remain3_2461);


wire[15:0] addr_selector3_2462;
wire[15:0] addr_remain3_2462;
address_decode_4 decoder_3_2462 = address_decode_4(addr_selector2_153[14],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2462,addr_remain3_2462);


wire[15:0] addr_selector3_2463;
wire[15:0] addr_remain3_2463;
address_decode_4 decoder_3_2463 = address_decode_4(addr_selector2_153[15],addr_remain2_153[15:0],addr_remain2_153,addr_selector3_2463,addr_remain3_2463);


wire[15:0] addr_selector3_2464;
wire[15:0] addr_remain3_2464;
address_decode_4 decoder_3_2464 = address_decode_4(addr_selector2_154[0],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2464,addr_remain3_2464);


wire[15:0] addr_selector3_2465;
wire[15:0] addr_remain3_2465;
address_decode_4 decoder_3_2465 = address_decode_4(addr_selector2_154[1],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2465,addr_remain3_2465);


wire[15:0] addr_selector3_2466;
wire[15:0] addr_remain3_2466;
address_decode_4 decoder_3_2466 = address_decode_4(addr_selector2_154[2],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2466,addr_remain3_2466);


wire[15:0] addr_selector3_2467;
wire[15:0] addr_remain3_2467;
address_decode_4 decoder_3_2467 = address_decode_4(addr_selector2_154[3],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2467,addr_remain3_2467);


wire[15:0] addr_selector3_2468;
wire[15:0] addr_remain3_2468;
address_decode_4 decoder_3_2468 = address_decode_4(addr_selector2_154[4],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2468,addr_remain3_2468);


wire[15:0] addr_selector3_2469;
wire[15:0] addr_remain3_2469;
address_decode_4 decoder_3_2469 = address_decode_4(addr_selector2_154[5],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2469,addr_remain3_2469);


wire[15:0] addr_selector3_2470;
wire[15:0] addr_remain3_2470;
address_decode_4 decoder_3_2470 = address_decode_4(addr_selector2_154[6],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2470,addr_remain3_2470);


wire[15:0] addr_selector3_2471;
wire[15:0] addr_remain3_2471;
address_decode_4 decoder_3_2471 = address_decode_4(addr_selector2_154[7],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2471,addr_remain3_2471);


wire[15:0] addr_selector3_2472;
wire[15:0] addr_remain3_2472;
address_decode_4 decoder_3_2472 = address_decode_4(addr_selector2_154[8],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2472,addr_remain3_2472);


wire[15:0] addr_selector3_2473;
wire[15:0] addr_remain3_2473;
address_decode_4 decoder_3_2473 = address_decode_4(addr_selector2_154[9],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2473,addr_remain3_2473);


wire[15:0] addr_selector3_2474;
wire[15:0] addr_remain3_2474;
address_decode_4 decoder_3_2474 = address_decode_4(addr_selector2_154[10],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2474,addr_remain3_2474);


wire[15:0] addr_selector3_2475;
wire[15:0] addr_remain3_2475;
address_decode_4 decoder_3_2475 = address_decode_4(addr_selector2_154[11],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2475,addr_remain3_2475);


wire[15:0] addr_selector3_2476;
wire[15:0] addr_remain3_2476;
address_decode_4 decoder_3_2476 = address_decode_4(addr_selector2_154[12],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2476,addr_remain3_2476);


wire[15:0] addr_selector3_2477;
wire[15:0] addr_remain3_2477;
address_decode_4 decoder_3_2477 = address_decode_4(addr_selector2_154[13],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2477,addr_remain3_2477);


wire[15:0] addr_selector3_2478;
wire[15:0] addr_remain3_2478;
address_decode_4 decoder_3_2478 = address_decode_4(addr_selector2_154[14],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2478,addr_remain3_2478);


wire[15:0] addr_selector3_2479;
wire[15:0] addr_remain3_2479;
address_decode_4 decoder_3_2479 = address_decode_4(addr_selector2_154[15],addr_remain2_154[15:0],addr_remain2_154,addr_selector3_2479,addr_remain3_2479);


wire[15:0] addr_selector3_2480;
wire[15:0] addr_remain3_2480;
address_decode_4 decoder_3_2480 = address_decode_4(addr_selector2_155[0],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2480,addr_remain3_2480);


wire[15:0] addr_selector3_2481;
wire[15:0] addr_remain3_2481;
address_decode_4 decoder_3_2481 = address_decode_4(addr_selector2_155[1],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2481,addr_remain3_2481);


wire[15:0] addr_selector3_2482;
wire[15:0] addr_remain3_2482;
address_decode_4 decoder_3_2482 = address_decode_4(addr_selector2_155[2],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2482,addr_remain3_2482);


wire[15:0] addr_selector3_2483;
wire[15:0] addr_remain3_2483;
address_decode_4 decoder_3_2483 = address_decode_4(addr_selector2_155[3],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2483,addr_remain3_2483);


wire[15:0] addr_selector3_2484;
wire[15:0] addr_remain3_2484;
address_decode_4 decoder_3_2484 = address_decode_4(addr_selector2_155[4],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2484,addr_remain3_2484);


wire[15:0] addr_selector3_2485;
wire[15:0] addr_remain3_2485;
address_decode_4 decoder_3_2485 = address_decode_4(addr_selector2_155[5],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2485,addr_remain3_2485);


wire[15:0] addr_selector3_2486;
wire[15:0] addr_remain3_2486;
address_decode_4 decoder_3_2486 = address_decode_4(addr_selector2_155[6],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2486,addr_remain3_2486);


wire[15:0] addr_selector3_2487;
wire[15:0] addr_remain3_2487;
address_decode_4 decoder_3_2487 = address_decode_4(addr_selector2_155[7],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2487,addr_remain3_2487);


wire[15:0] addr_selector3_2488;
wire[15:0] addr_remain3_2488;
address_decode_4 decoder_3_2488 = address_decode_4(addr_selector2_155[8],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2488,addr_remain3_2488);


wire[15:0] addr_selector3_2489;
wire[15:0] addr_remain3_2489;
address_decode_4 decoder_3_2489 = address_decode_4(addr_selector2_155[9],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2489,addr_remain3_2489);


wire[15:0] addr_selector3_2490;
wire[15:0] addr_remain3_2490;
address_decode_4 decoder_3_2490 = address_decode_4(addr_selector2_155[10],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2490,addr_remain3_2490);


wire[15:0] addr_selector3_2491;
wire[15:0] addr_remain3_2491;
address_decode_4 decoder_3_2491 = address_decode_4(addr_selector2_155[11],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2491,addr_remain3_2491);


wire[15:0] addr_selector3_2492;
wire[15:0] addr_remain3_2492;
address_decode_4 decoder_3_2492 = address_decode_4(addr_selector2_155[12],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2492,addr_remain3_2492);


wire[15:0] addr_selector3_2493;
wire[15:0] addr_remain3_2493;
address_decode_4 decoder_3_2493 = address_decode_4(addr_selector2_155[13],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2493,addr_remain3_2493);


wire[15:0] addr_selector3_2494;
wire[15:0] addr_remain3_2494;
address_decode_4 decoder_3_2494 = address_decode_4(addr_selector2_155[14],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2494,addr_remain3_2494);


wire[15:0] addr_selector3_2495;
wire[15:0] addr_remain3_2495;
address_decode_4 decoder_3_2495 = address_decode_4(addr_selector2_155[15],addr_remain2_155[15:0],addr_remain2_155,addr_selector3_2495,addr_remain3_2495);


wire[15:0] addr_selector3_2496;
wire[15:0] addr_remain3_2496;
address_decode_4 decoder_3_2496 = address_decode_4(addr_selector2_156[0],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2496,addr_remain3_2496);


wire[15:0] addr_selector3_2497;
wire[15:0] addr_remain3_2497;
address_decode_4 decoder_3_2497 = address_decode_4(addr_selector2_156[1],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2497,addr_remain3_2497);


wire[15:0] addr_selector3_2498;
wire[15:0] addr_remain3_2498;
address_decode_4 decoder_3_2498 = address_decode_4(addr_selector2_156[2],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2498,addr_remain3_2498);


wire[15:0] addr_selector3_2499;
wire[15:0] addr_remain3_2499;
address_decode_4 decoder_3_2499 = address_decode_4(addr_selector2_156[3],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2499,addr_remain3_2499);


wire[15:0] addr_selector3_2500;
wire[15:0] addr_remain3_2500;
address_decode_4 decoder_3_2500 = address_decode_4(addr_selector2_156[4],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2500,addr_remain3_2500);


wire[15:0] addr_selector3_2501;
wire[15:0] addr_remain3_2501;
address_decode_4 decoder_3_2501 = address_decode_4(addr_selector2_156[5],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2501,addr_remain3_2501);


wire[15:0] addr_selector3_2502;
wire[15:0] addr_remain3_2502;
address_decode_4 decoder_3_2502 = address_decode_4(addr_selector2_156[6],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2502,addr_remain3_2502);


wire[15:0] addr_selector3_2503;
wire[15:0] addr_remain3_2503;
address_decode_4 decoder_3_2503 = address_decode_4(addr_selector2_156[7],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2503,addr_remain3_2503);


wire[15:0] addr_selector3_2504;
wire[15:0] addr_remain3_2504;
address_decode_4 decoder_3_2504 = address_decode_4(addr_selector2_156[8],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2504,addr_remain3_2504);


wire[15:0] addr_selector3_2505;
wire[15:0] addr_remain3_2505;
address_decode_4 decoder_3_2505 = address_decode_4(addr_selector2_156[9],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2505,addr_remain3_2505);


wire[15:0] addr_selector3_2506;
wire[15:0] addr_remain3_2506;
address_decode_4 decoder_3_2506 = address_decode_4(addr_selector2_156[10],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2506,addr_remain3_2506);


wire[15:0] addr_selector3_2507;
wire[15:0] addr_remain3_2507;
address_decode_4 decoder_3_2507 = address_decode_4(addr_selector2_156[11],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2507,addr_remain3_2507);


wire[15:0] addr_selector3_2508;
wire[15:0] addr_remain3_2508;
address_decode_4 decoder_3_2508 = address_decode_4(addr_selector2_156[12],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2508,addr_remain3_2508);


wire[15:0] addr_selector3_2509;
wire[15:0] addr_remain3_2509;
address_decode_4 decoder_3_2509 = address_decode_4(addr_selector2_156[13],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2509,addr_remain3_2509);


wire[15:0] addr_selector3_2510;
wire[15:0] addr_remain3_2510;
address_decode_4 decoder_3_2510 = address_decode_4(addr_selector2_156[14],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2510,addr_remain3_2510);


wire[15:0] addr_selector3_2511;
wire[15:0] addr_remain3_2511;
address_decode_4 decoder_3_2511 = address_decode_4(addr_selector2_156[15],addr_remain2_156[15:0],addr_remain2_156,addr_selector3_2511,addr_remain3_2511);


wire[15:0] addr_selector3_2512;
wire[15:0] addr_remain3_2512;
address_decode_4 decoder_3_2512 = address_decode_4(addr_selector2_157[0],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2512,addr_remain3_2512);


wire[15:0] addr_selector3_2513;
wire[15:0] addr_remain3_2513;
address_decode_4 decoder_3_2513 = address_decode_4(addr_selector2_157[1],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2513,addr_remain3_2513);


wire[15:0] addr_selector3_2514;
wire[15:0] addr_remain3_2514;
address_decode_4 decoder_3_2514 = address_decode_4(addr_selector2_157[2],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2514,addr_remain3_2514);


wire[15:0] addr_selector3_2515;
wire[15:0] addr_remain3_2515;
address_decode_4 decoder_3_2515 = address_decode_4(addr_selector2_157[3],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2515,addr_remain3_2515);


wire[15:0] addr_selector3_2516;
wire[15:0] addr_remain3_2516;
address_decode_4 decoder_3_2516 = address_decode_4(addr_selector2_157[4],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2516,addr_remain3_2516);


wire[15:0] addr_selector3_2517;
wire[15:0] addr_remain3_2517;
address_decode_4 decoder_3_2517 = address_decode_4(addr_selector2_157[5],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2517,addr_remain3_2517);


wire[15:0] addr_selector3_2518;
wire[15:0] addr_remain3_2518;
address_decode_4 decoder_3_2518 = address_decode_4(addr_selector2_157[6],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2518,addr_remain3_2518);


wire[15:0] addr_selector3_2519;
wire[15:0] addr_remain3_2519;
address_decode_4 decoder_3_2519 = address_decode_4(addr_selector2_157[7],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2519,addr_remain3_2519);


wire[15:0] addr_selector3_2520;
wire[15:0] addr_remain3_2520;
address_decode_4 decoder_3_2520 = address_decode_4(addr_selector2_157[8],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2520,addr_remain3_2520);


wire[15:0] addr_selector3_2521;
wire[15:0] addr_remain3_2521;
address_decode_4 decoder_3_2521 = address_decode_4(addr_selector2_157[9],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2521,addr_remain3_2521);


wire[15:0] addr_selector3_2522;
wire[15:0] addr_remain3_2522;
address_decode_4 decoder_3_2522 = address_decode_4(addr_selector2_157[10],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2522,addr_remain3_2522);


wire[15:0] addr_selector3_2523;
wire[15:0] addr_remain3_2523;
address_decode_4 decoder_3_2523 = address_decode_4(addr_selector2_157[11],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2523,addr_remain3_2523);


wire[15:0] addr_selector3_2524;
wire[15:0] addr_remain3_2524;
address_decode_4 decoder_3_2524 = address_decode_4(addr_selector2_157[12],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2524,addr_remain3_2524);


wire[15:0] addr_selector3_2525;
wire[15:0] addr_remain3_2525;
address_decode_4 decoder_3_2525 = address_decode_4(addr_selector2_157[13],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2525,addr_remain3_2525);


wire[15:0] addr_selector3_2526;
wire[15:0] addr_remain3_2526;
address_decode_4 decoder_3_2526 = address_decode_4(addr_selector2_157[14],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2526,addr_remain3_2526);


wire[15:0] addr_selector3_2527;
wire[15:0] addr_remain3_2527;
address_decode_4 decoder_3_2527 = address_decode_4(addr_selector2_157[15],addr_remain2_157[15:0],addr_remain2_157,addr_selector3_2527,addr_remain3_2527);


wire[15:0] addr_selector3_2528;
wire[15:0] addr_remain3_2528;
address_decode_4 decoder_3_2528 = address_decode_4(addr_selector2_158[0],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2528,addr_remain3_2528);


wire[15:0] addr_selector3_2529;
wire[15:0] addr_remain3_2529;
address_decode_4 decoder_3_2529 = address_decode_4(addr_selector2_158[1],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2529,addr_remain3_2529);


wire[15:0] addr_selector3_2530;
wire[15:0] addr_remain3_2530;
address_decode_4 decoder_3_2530 = address_decode_4(addr_selector2_158[2],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2530,addr_remain3_2530);


wire[15:0] addr_selector3_2531;
wire[15:0] addr_remain3_2531;
address_decode_4 decoder_3_2531 = address_decode_4(addr_selector2_158[3],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2531,addr_remain3_2531);


wire[15:0] addr_selector3_2532;
wire[15:0] addr_remain3_2532;
address_decode_4 decoder_3_2532 = address_decode_4(addr_selector2_158[4],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2532,addr_remain3_2532);


wire[15:0] addr_selector3_2533;
wire[15:0] addr_remain3_2533;
address_decode_4 decoder_3_2533 = address_decode_4(addr_selector2_158[5],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2533,addr_remain3_2533);


wire[15:0] addr_selector3_2534;
wire[15:0] addr_remain3_2534;
address_decode_4 decoder_3_2534 = address_decode_4(addr_selector2_158[6],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2534,addr_remain3_2534);


wire[15:0] addr_selector3_2535;
wire[15:0] addr_remain3_2535;
address_decode_4 decoder_3_2535 = address_decode_4(addr_selector2_158[7],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2535,addr_remain3_2535);


wire[15:0] addr_selector3_2536;
wire[15:0] addr_remain3_2536;
address_decode_4 decoder_3_2536 = address_decode_4(addr_selector2_158[8],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2536,addr_remain3_2536);


wire[15:0] addr_selector3_2537;
wire[15:0] addr_remain3_2537;
address_decode_4 decoder_3_2537 = address_decode_4(addr_selector2_158[9],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2537,addr_remain3_2537);


wire[15:0] addr_selector3_2538;
wire[15:0] addr_remain3_2538;
address_decode_4 decoder_3_2538 = address_decode_4(addr_selector2_158[10],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2538,addr_remain3_2538);


wire[15:0] addr_selector3_2539;
wire[15:0] addr_remain3_2539;
address_decode_4 decoder_3_2539 = address_decode_4(addr_selector2_158[11],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2539,addr_remain3_2539);


wire[15:0] addr_selector3_2540;
wire[15:0] addr_remain3_2540;
address_decode_4 decoder_3_2540 = address_decode_4(addr_selector2_158[12],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2540,addr_remain3_2540);


wire[15:0] addr_selector3_2541;
wire[15:0] addr_remain3_2541;
address_decode_4 decoder_3_2541 = address_decode_4(addr_selector2_158[13],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2541,addr_remain3_2541);


wire[15:0] addr_selector3_2542;
wire[15:0] addr_remain3_2542;
address_decode_4 decoder_3_2542 = address_decode_4(addr_selector2_158[14],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2542,addr_remain3_2542);


wire[15:0] addr_selector3_2543;
wire[15:0] addr_remain3_2543;
address_decode_4 decoder_3_2543 = address_decode_4(addr_selector2_158[15],addr_remain2_158[15:0],addr_remain2_158,addr_selector3_2543,addr_remain3_2543);


wire[15:0] addr_selector3_2544;
wire[15:0] addr_remain3_2544;
address_decode_4 decoder_3_2544 = address_decode_4(addr_selector2_159[0],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2544,addr_remain3_2544);


wire[15:0] addr_selector3_2545;
wire[15:0] addr_remain3_2545;
address_decode_4 decoder_3_2545 = address_decode_4(addr_selector2_159[1],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2545,addr_remain3_2545);


wire[15:0] addr_selector3_2546;
wire[15:0] addr_remain3_2546;
address_decode_4 decoder_3_2546 = address_decode_4(addr_selector2_159[2],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2546,addr_remain3_2546);


wire[15:0] addr_selector3_2547;
wire[15:0] addr_remain3_2547;
address_decode_4 decoder_3_2547 = address_decode_4(addr_selector2_159[3],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2547,addr_remain3_2547);


wire[15:0] addr_selector3_2548;
wire[15:0] addr_remain3_2548;
address_decode_4 decoder_3_2548 = address_decode_4(addr_selector2_159[4],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2548,addr_remain3_2548);


wire[15:0] addr_selector3_2549;
wire[15:0] addr_remain3_2549;
address_decode_4 decoder_3_2549 = address_decode_4(addr_selector2_159[5],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2549,addr_remain3_2549);


wire[15:0] addr_selector3_2550;
wire[15:0] addr_remain3_2550;
address_decode_4 decoder_3_2550 = address_decode_4(addr_selector2_159[6],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2550,addr_remain3_2550);


wire[15:0] addr_selector3_2551;
wire[15:0] addr_remain3_2551;
address_decode_4 decoder_3_2551 = address_decode_4(addr_selector2_159[7],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2551,addr_remain3_2551);


wire[15:0] addr_selector3_2552;
wire[15:0] addr_remain3_2552;
address_decode_4 decoder_3_2552 = address_decode_4(addr_selector2_159[8],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2552,addr_remain3_2552);


wire[15:0] addr_selector3_2553;
wire[15:0] addr_remain3_2553;
address_decode_4 decoder_3_2553 = address_decode_4(addr_selector2_159[9],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2553,addr_remain3_2553);


wire[15:0] addr_selector3_2554;
wire[15:0] addr_remain3_2554;
address_decode_4 decoder_3_2554 = address_decode_4(addr_selector2_159[10],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2554,addr_remain3_2554);


wire[15:0] addr_selector3_2555;
wire[15:0] addr_remain3_2555;
address_decode_4 decoder_3_2555 = address_decode_4(addr_selector2_159[11],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2555,addr_remain3_2555);


wire[15:0] addr_selector3_2556;
wire[15:0] addr_remain3_2556;
address_decode_4 decoder_3_2556 = address_decode_4(addr_selector2_159[12],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2556,addr_remain3_2556);


wire[15:0] addr_selector3_2557;
wire[15:0] addr_remain3_2557;
address_decode_4 decoder_3_2557 = address_decode_4(addr_selector2_159[13],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2557,addr_remain3_2557);


wire[15:0] addr_selector3_2558;
wire[15:0] addr_remain3_2558;
address_decode_4 decoder_3_2558 = address_decode_4(addr_selector2_159[14],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2558,addr_remain3_2558);


wire[15:0] addr_selector3_2559;
wire[15:0] addr_remain3_2559;
address_decode_4 decoder_3_2559 = address_decode_4(addr_selector2_159[15],addr_remain2_159[15:0],addr_remain2_159,addr_selector3_2559,addr_remain3_2559);


wire[15:0] addr_selector3_2560;
wire[15:0] addr_remain3_2560;
address_decode_4 decoder_3_2560 = address_decode_4(addr_selector2_160[0],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2560,addr_remain3_2560);


wire[15:0] addr_selector3_2561;
wire[15:0] addr_remain3_2561;
address_decode_4 decoder_3_2561 = address_decode_4(addr_selector2_160[1],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2561,addr_remain3_2561);


wire[15:0] addr_selector3_2562;
wire[15:0] addr_remain3_2562;
address_decode_4 decoder_3_2562 = address_decode_4(addr_selector2_160[2],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2562,addr_remain3_2562);


wire[15:0] addr_selector3_2563;
wire[15:0] addr_remain3_2563;
address_decode_4 decoder_3_2563 = address_decode_4(addr_selector2_160[3],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2563,addr_remain3_2563);


wire[15:0] addr_selector3_2564;
wire[15:0] addr_remain3_2564;
address_decode_4 decoder_3_2564 = address_decode_4(addr_selector2_160[4],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2564,addr_remain3_2564);


wire[15:0] addr_selector3_2565;
wire[15:0] addr_remain3_2565;
address_decode_4 decoder_3_2565 = address_decode_4(addr_selector2_160[5],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2565,addr_remain3_2565);


wire[15:0] addr_selector3_2566;
wire[15:0] addr_remain3_2566;
address_decode_4 decoder_3_2566 = address_decode_4(addr_selector2_160[6],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2566,addr_remain3_2566);


wire[15:0] addr_selector3_2567;
wire[15:0] addr_remain3_2567;
address_decode_4 decoder_3_2567 = address_decode_4(addr_selector2_160[7],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2567,addr_remain3_2567);


wire[15:0] addr_selector3_2568;
wire[15:0] addr_remain3_2568;
address_decode_4 decoder_3_2568 = address_decode_4(addr_selector2_160[8],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2568,addr_remain3_2568);


wire[15:0] addr_selector3_2569;
wire[15:0] addr_remain3_2569;
address_decode_4 decoder_3_2569 = address_decode_4(addr_selector2_160[9],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2569,addr_remain3_2569);


wire[15:0] addr_selector3_2570;
wire[15:0] addr_remain3_2570;
address_decode_4 decoder_3_2570 = address_decode_4(addr_selector2_160[10],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2570,addr_remain3_2570);


wire[15:0] addr_selector3_2571;
wire[15:0] addr_remain3_2571;
address_decode_4 decoder_3_2571 = address_decode_4(addr_selector2_160[11],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2571,addr_remain3_2571);


wire[15:0] addr_selector3_2572;
wire[15:0] addr_remain3_2572;
address_decode_4 decoder_3_2572 = address_decode_4(addr_selector2_160[12],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2572,addr_remain3_2572);


wire[15:0] addr_selector3_2573;
wire[15:0] addr_remain3_2573;
address_decode_4 decoder_3_2573 = address_decode_4(addr_selector2_160[13],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2573,addr_remain3_2573);


wire[15:0] addr_selector3_2574;
wire[15:0] addr_remain3_2574;
address_decode_4 decoder_3_2574 = address_decode_4(addr_selector2_160[14],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2574,addr_remain3_2574);


wire[15:0] addr_selector3_2575;
wire[15:0] addr_remain3_2575;
address_decode_4 decoder_3_2575 = address_decode_4(addr_selector2_160[15],addr_remain2_160[15:0],addr_remain2_160,addr_selector3_2575,addr_remain3_2575);


wire[15:0] addr_selector3_2576;
wire[15:0] addr_remain3_2576;
address_decode_4 decoder_3_2576 = address_decode_4(addr_selector2_161[0],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2576,addr_remain3_2576);


wire[15:0] addr_selector3_2577;
wire[15:0] addr_remain3_2577;
address_decode_4 decoder_3_2577 = address_decode_4(addr_selector2_161[1],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2577,addr_remain3_2577);


wire[15:0] addr_selector3_2578;
wire[15:0] addr_remain3_2578;
address_decode_4 decoder_3_2578 = address_decode_4(addr_selector2_161[2],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2578,addr_remain3_2578);


wire[15:0] addr_selector3_2579;
wire[15:0] addr_remain3_2579;
address_decode_4 decoder_3_2579 = address_decode_4(addr_selector2_161[3],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2579,addr_remain3_2579);


wire[15:0] addr_selector3_2580;
wire[15:0] addr_remain3_2580;
address_decode_4 decoder_3_2580 = address_decode_4(addr_selector2_161[4],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2580,addr_remain3_2580);


wire[15:0] addr_selector3_2581;
wire[15:0] addr_remain3_2581;
address_decode_4 decoder_3_2581 = address_decode_4(addr_selector2_161[5],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2581,addr_remain3_2581);


wire[15:0] addr_selector3_2582;
wire[15:0] addr_remain3_2582;
address_decode_4 decoder_3_2582 = address_decode_4(addr_selector2_161[6],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2582,addr_remain3_2582);


wire[15:0] addr_selector3_2583;
wire[15:0] addr_remain3_2583;
address_decode_4 decoder_3_2583 = address_decode_4(addr_selector2_161[7],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2583,addr_remain3_2583);


wire[15:0] addr_selector3_2584;
wire[15:0] addr_remain3_2584;
address_decode_4 decoder_3_2584 = address_decode_4(addr_selector2_161[8],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2584,addr_remain3_2584);


wire[15:0] addr_selector3_2585;
wire[15:0] addr_remain3_2585;
address_decode_4 decoder_3_2585 = address_decode_4(addr_selector2_161[9],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2585,addr_remain3_2585);


wire[15:0] addr_selector3_2586;
wire[15:0] addr_remain3_2586;
address_decode_4 decoder_3_2586 = address_decode_4(addr_selector2_161[10],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2586,addr_remain3_2586);


wire[15:0] addr_selector3_2587;
wire[15:0] addr_remain3_2587;
address_decode_4 decoder_3_2587 = address_decode_4(addr_selector2_161[11],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2587,addr_remain3_2587);


wire[15:0] addr_selector3_2588;
wire[15:0] addr_remain3_2588;
address_decode_4 decoder_3_2588 = address_decode_4(addr_selector2_161[12],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2588,addr_remain3_2588);


wire[15:0] addr_selector3_2589;
wire[15:0] addr_remain3_2589;
address_decode_4 decoder_3_2589 = address_decode_4(addr_selector2_161[13],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2589,addr_remain3_2589);


wire[15:0] addr_selector3_2590;
wire[15:0] addr_remain3_2590;
address_decode_4 decoder_3_2590 = address_decode_4(addr_selector2_161[14],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2590,addr_remain3_2590);


wire[15:0] addr_selector3_2591;
wire[15:0] addr_remain3_2591;
address_decode_4 decoder_3_2591 = address_decode_4(addr_selector2_161[15],addr_remain2_161[15:0],addr_remain2_161,addr_selector3_2591,addr_remain3_2591);


wire[15:0] addr_selector3_2592;
wire[15:0] addr_remain3_2592;
address_decode_4 decoder_3_2592 = address_decode_4(addr_selector2_162[0],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2592,addr_remain3_2592);


wire[15:0] addr_selector3_2593;
wire[15:0] addr_remain3_2593;
address_decode_4 decoder_3_2593 = address_decode_4(addr_selector2_162[1],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2593,addr_remain3_2593);


wire[15:0] addr_selector3_2594;
wire[15:0] addr_remain3_2594;
address_decode_4 decoder_3_2594 = address_decode_4(addr_selector2_162[2],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2594,addr_remain3_2594);


wire[15:0] addr_selector3_2595;
wire[15:0] addr_remain3_2595;
address_decode_4 decoder_3_2595 = address_decode_4(addr_selector2_162[3],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2595,addr_remain3_2595);


wire[15:0] addr_selector3_2596;
wire[15:0] addr_remain3_2596;
address_decode_4 decoder_3_2596 = address_decode_4(addr_selector2_162[4],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2596,addr_remain3_2596);


wire[15:0] addr_selector3_2597;
wire[15:0] addr_remain3_2597;
address_decode_4 decoder_3_2597 = address_decode_4(addr_selector2_162[5],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2597,addr_remain3_2597);


wire[15:0] addr_selector3_2598;
wire[15:0] addr_remain3_2598;
address_decode_4 decoder_3_2598 = address_decode_4(addr_selector2_162[6],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2598,addr_remain3_2598);


wire[15:0] addr_selector3_2599;
wire[15:0] addr_remain3_2599;
address_decode_4 decoder_3_2599 = address_decode_4(addr_selector2_162[7],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2599,addr_remain3_2599);


wire[15:0] addr_selector3_2600;
wire[15:0] addr_remain3_2600;
address_decode_4 decoder_3_2600 = address_decode_4(addr_selector2_162[8],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2600,addr_remain3_2600);


wire[15:0] addr_selector3_2601;
wire[15:0] addr_remain3_2601;
address_decode_4 decoder_3_2601 = address_decode_4(addr_selector2_162[9],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2601,addr_remain3_2601);


wire[15:0] addr_selector3_2602;
wire[15:0] addr_remain3_2602;
address_decode_4 decoder_3_2602 = address_decode_4(addr_selector2_162[10],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2602,addr_remain3_2602);


wire[15:0] addr_selector3_2603;
wire[15:0] addr_remain3_2603;
address_decode_4 decoder_3_2603 = address_decode_4(addr_selector2_162[11],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2603,addr_remain3_2603);


wire[15:0] addr_selector3_2604;
wire[15:0] addr_remain3_2604;
address_decode_4 decoder_3_2604 = address_decode_4(addr_selector2_162[12],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2604,addr_remain3_2604);


wire[15:0] addr_selector3_2605;
wire[15:0] addr_remain3_2605;
address_decode_4 decoder_3_2605 = address_decode_4(addr_selector2_162[13],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2605,addr_remain3_2605);


wire[15:0] addr_selector3_2606;
wire[15:0] addr_remain3_2606;
address_decode_4 decoder_3_2606 = address_decode_4(addr_selector2_162[14],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2606,addr_remain3_2606);


wire[15:0] addr_selector3_2607;
wire[15:0] addr_remain3_2607;
address_decode_4 decoder_3_2607 = address_decode_4(addr_selector2_162[15],addr_remain2_162[15:0],addr_remain2_162,addr_selector3_2607,addr_remain3_2607);


wire[15:0] addr_selector3_2608;
wire[15:0] addr_remain3_2608;
address_decode_4 decoder_3_2608 = address_decode_4(addr_selector2_163[0],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2608,addr_remain3_2608);


wire[15:0] addr_selector3_2609;
wire[15:0] addr_remain3_2609;
address_decode_4 decoder_3_2609 = address_decode_4(addr_selector2_163[1],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2609,addr_remain3_2609);


wire[15:0] addr_selector3_2610;
wire[15:0] addr_remain3_2610;
address_decode_4 decoder_3_2610 = address_decode_4(addr_selector2_163[2],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2610,addr_remain3_2610);


wire[15:0] addr_selector3_2611;
wire[15:0] addr_remain3_2611;
address_decode_4 decoder_3_2611 = address_decode_4(addr_selector2_163[3],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2611,addr_remain3_2611);


wire[15:0] addr_selector3_2612;
wire[15:0] addr_remain3_2612;
address_decode_4 decoder_3_2612 = address_decode_4(addr_selector2_163[4],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2612,addr_remain3_2612);


wire[15:0] addr_selector3_2613;
wire[15:0] addr_remain3_2613;
address_decode_4 decoder_3_2613 = address_decode_4(addr_selector2_163[5],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2613,addr_remain3_2613);


wire[15:0] addr_selector3_2614;
wire[15:0] addr_remain3_2614;
address_decode_4 decoder_3_2614 = address_decode_4(addr_selector2_163[6],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2614,addr_remain3_2614);


wire[15:0] addr_selector3_2615;
wire[15:0] addr_remain3_2615;
address_decode_4 decoder_3_2615 = address_decode_4(addr_selector2_163[7],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2615,addr_remain3_2615);


wire[15:0] addr_selector3_2616;
wire[15:0] addr_remain3_2616;
address_decode_4 decoder_3_2616 = address_decode_4(addr_selector2_163[8],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2616,addr_remain3_2616);


wire[15:0] addr_selector3_2617;
wire[15:0] addr_remain3_2617;
address_decode_4 decoder_3_2617 = address_decode_4(addr_selector2_163[9],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2617,addr_remain3_2617);


wire[15:0] addr_selector3_2618;
wire[15:0] addr_remain3_2618;
address_decode_4 decoder_3_2618 = address_decode_4(addr_selector2_163[10],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2618,addr_remain3_2618);


wire[15:0] addr_selector3_2619;
wire[15:0] addr_remain3_2619;
address_decode_4 decoder_3_2619 = address_decode_4(addr_selector2_163[11],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2619,addr_remain3_2619);


wire[15:0] addr_selector3_2620;
wire[15:0] addr_remain3_2620;
address_decode_4 decoder_3_2620 = address_decode_4(addr_selector2_163[12],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2620,addr_remain3_2620);


wire[15:0] addr_selector3_2621;
wire[15:0] addr_remain3_2621;
address_decode_4 decoder_3_2621 = address_decode_4(addr_selector2_163[13],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2621,addr_remain3_2621);


wire[15:0] addr_selector3_2622;
wire[15:0] addr_remain3_2622;
address_decode_4 decoder_3_2622 = address_decode_4(addr_selector2_163[14],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2622,addr_remain3_2622);


wire[15:0] addr_selector3_2623;
wire[15:0] addr_remain3_2623;
address_decode_4 decoder_3_2623 = address_decode_4(addr_selector2_163[15],addr_remain2_163[15:0],addr_remain2_163,addr_selector3_2623,addr_remain3_2623);


wire[15:0] addr_selector3_2624;
wire[15:0] addr_remain3_2624;
address_decode_4 decoder_3_2624 = address_decode_4(addr_selector2_164[0],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2624,addr_remain3_2624);


wire[15:0] addr_selector3_2625;
wire[15:0] addr_remain3_2625;
address_decode_4 decoder_3_2625 = address_decode_4(addr_selector2_164[1],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2625,addr_remain3_2625);


wire[15:0] addr_selector3_2626;
wire[15:0] addr_remain3_2626;
address_decode_4 decoder_3_2626 = address_decode_4(addr_selector2_164[2],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2626,addr_remain3_2626);


wire[15:0] addr_selector3_2627;
wire[15:0] addr_remain3_2627;
address_decode_4 decoder_3_2627 = address_decode_4(addr_selector2_164[3],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2627,addr_remain3_2627);


wire[15:0] addr_selector3_2628;
wire[15:0] addr_remain3_2628;
address_decode_4 decoder_3_2628 = address_decode_4(addr_selector2_164[4],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2628,addr_remain3_2628);


wire[15:0] addr_selector3_2629;
wire[15:0] addr_remain3_2629;
address_decode_4 decoder_3_2629 = address_decode_4(addr_selector2_164[5],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2629,addr_remain3_2629);


wire[15:0] addr_selector3_2630;
wire[15:0] addr_remain3_2630;
address_decode_4 decoder_3_2630 = address_decode_4(addr_selector2_164[6],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2630,addr_remain3_2630);


wire[15:0] addr_selector3_2631;
wire[15:0] addr_remain3_2631;
address_decode_4 decoder_3_2631 = address_decode_4(addr_selector2_164[7],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2631,addr_remain3_2631);


wire[15:0] addr_selector3_2632;
wire[15:0] addr_remain3_2632;
address_decode_4 decoder_3_2632 = address_decode_4(addr_selector2_164[8],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2632,addr_remain3_2632);


wire[15:0] addr_selector3_2633;
wire[15:0] addr_remain3_2633;
address_decode_4 decoder_3_2633 = address_decode_4(addr_selector2_164[9],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2633,addr_remain3_2633);


wire[15:0] addr_selector3_2634;
wire[15:0] addr_remain3_2634;
address_decode_4 decoder_3_2634 = address_decode_4(addr_selector2_164[10],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2634,addr_remain3_2634);


wire[15:0] addr_selector3_2635;
wire[15:0] addr_remain3_2635;
address_decode_4 decoder_3_2635 = address_decode_4(addr_selector2_164[11],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2635,addr_remain3_2635);


wire[15:0] addr_selector3_2636;
wire[15:0] addr_remain3_2636;
address_decode_4 decoder_3_2636 = address_decode_4(addr_selector2_164[12],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2636,addr_remain3_2636);


wire[15:0] addr_selector3_2637;
wire[15:0] addr_remain3_2637;
address_decode_4 decoder_3_2637 = address_decode_4(addr_selector2_164[13],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2637,addr_remain3_2637);


wire[15:0] addr_selector3_2638;
wire[15:0] addr_remain3_2638;
address_decode_4 decoder_3_2638 = address_decode_4(addr_selector2_164[14],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2638,addr_remain3_2638);


wire[15:0] addr_selector3_2639;
wire[15:0] addr_remain3_2639;
address_decode_4 decoder_3_2639 = address_decode_4(addr_selector2_164[15],addr_remain2_164[15:0],addr_remain2_164,addr_selector3_2639,addr_remain3_2639);


wire[15:0] addr_selector3_2640;
wire[15:0] addr_remain3_2640;
address_decode_4 decoder_3_2640 = address_decode_4(addr_selector2_165[0],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2640,addr_remain3_2640);


wire[15:0] addr_selector3_2641;
wire[15:0] addr_remain3_2641;
address_decode_4 decoder_3_2641 = address_decode_4(addr_selector2_165[1],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2641,addr_remain3_2641);


wire[15:0] addr_selector3_2642;
wire[15:0] addr_remain3_2642;
address_decode_4 decoder_3_2642 = address_decode_4(addr_selector2_165[2],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2642,addr_remain3_2642);


wire[15:0] addr_selector3_2643;
wire[15:0] addr_remain3_2643;
address_decode_4 decoder_3_2643 = address_decode_4(addr_selector2_165[3],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2643,addr_remain3_2643);


wire[15:0] addr_selector3_2644;
wire[15:0] addr_remain3_2644;
address_decode_4 decoder_3_2644 = address_decode_4(addr_selector2_165[4],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2644,addr_remain3_2644);


wire[15:0] addr_selector3_2645;
wire[15:0] addr_remain3_2645;
address_decode_4 decoder_3_2645 = address_decode_4(addr_selector2_165[5],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2645,addr_remain3_2645);


wire[15:0] addr_selector3_2646;
wire[15:0] addr_remain3_2646;
address_decode_4 decoder_3_2646 = address_decode_4(addr_selector2_165[6],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2646,addr_remain3_2646);


wire[15:0] addr_selector3_2647;
wire[15:0] addr_remain3_2647;
address_decode_4 decoder_3_2647 = address_decode_4(addr_selector2_165[7],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2647,addr_remain3_2647);


wire[15:0] addr_selector3_2648;
wire[15:0] addr_remain3_2648;
address_decode_4 decoder_3_2648 = address_decode_4(addr_selector2_165[8],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2648,addr_remain3_2648);


wire[15:0] addr_selector3_2649;
wire[15:0] addr_remain3_2649;
address_decode_4 decoder_3_2649 = address_decode_4(addr_selector2_165[9],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2649,addr_remain3_2649);


wire[15:0] addr_selector3_2650;
wire[15:0] addr_remain3_2650;
address_decode_4 decoder_3_2650 = address_decode_4(addr_selector2_165[10],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2650,addr_remain3_2650);


wire[15:0] addr_selector3_2651;
wire[15:0] addr_remain3_2651;
address_decode_4 decoder_3_2651 = address_decode_4(addr_selector2_165[11],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2651,addr_remain3_2651);


wire[15:0] addr_selector3_2652;
wire[15:0] addr_remain3_2652;
address_decode_4 decoder_3_2652 = address_decode_4(addr_selector2_165[12],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2652,addr_remain3_2652);


wire[15:0] addr_selector3_2653;
wire[15:0] addr_remain3_2653;
address_decode_4 decoder_3_2653 = address_decode_4(addr_selector2_165[13],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2653,addr_remain3_2653);


wire[15:0] addr_selector3_2654;
wire[15:0] addr_remain3_2654;
address_decode_4 decoder_3_2654 = address_decode_4(addr_selector2_165[14],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2654,addr_remain3_2654);


wire[15:0] addr_selector3_2655;
wire[15:0] addr_remain3_2655;
address_decode_4 decoder_3_2655 = address_decode_4(addr_selector2_165[15],addr_remain2_165[15:0],addr_remain2_165,addr_selector3_2655,addr_remain3_2655);


wire[15:0] addr_selector3_2656;
wire[15:0] addr_remain3_2656;
address_decode_4 decoder_3_2656 = address_decode_4(addr_selector2_166[0],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2656,addr_remain3_2656);


wire[15:0] addr_selector3_2657;
wire[15:0] addr_remain3_2657;
address_decode_4 decoder_3_2657 = address_decode_4(addr_selector2_166[1],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2657,addr_remain3_2657);


wire[15:0] addr_selector3_2658;
wire[15:0] addr_remain3_2658;
address_decode_4 decoder_3_2658 = address_decode_4(addr_selector2_166[2],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2658,addr_remain3_2658);


wire[15:0] addr_selector3_2659;
wire[15:0] addr_remain3_2659;
address_decode_4 decoder_3_2659 = address_decode_4(addr_selector2_166[3],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2659,addr_remain3_2659);


wire[15:0] addr_selector3_2660;
wire[15:0] addr_remain3_2660;
address_decode_4 decoder_3_2660 = address_decode_4(addr_selector2_166[4],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2660,addr_remain3_2660);


wire[15:0] addr_selector3_2661;
wire[15:0] addr_remain3_2661;
address_decode_4 decoder_3_2661 = address_decode_4(addr_selector2_166[5],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2661,addr_remain3_2661);


wire[15:0] addr_selector3_2662;
wire[15:0] addr_remain3_2662;
address_decode_4 decoder_3_2662 = address_decode_4(addr_selector2_166[6],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2662,addr_remain3_2662);


wire[15:0] addr_selector3_2663;
wire[15:0] addr_remain3_2663;
address_decode_4 decoder_3_2663 = address_decode_4(addr_selector2_166[7],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2663,addr_remain3_2663);


wire[15:0] addr_selector3_2664;
wire[15:0] addr_remain3_2664;
address_decode_4 decoder_3_2664 = address_decode_4(addr_selector2_166[8],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2664,addr_remain3_2664);


wire[15:0] addr_selector3_2665;
wire[15:0] addr_remain3_2665;
address_decode_4 decoder_3_2665 = address_decode_4(addr_selector2_166[9],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2665,addr_remain3_2665);


wire[15:0] addr_selector3_2666;
wire[15:0] addr_remain3_2666;
address_decode_4 decoder_3_2666 = address_decode_4(addr_selector2_166[10],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2666,addr_remain3_2666);


wire[15:0] addr_selector3_2667;
wire[15:0] addr_remain3_2667;
address_decode_4 decoder_3_2667 = address_decode_4(addr_selector2_166[11],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2667,addr_remain3_2667);


wire[15:0] addr_selector3_2668;
wire[15:0] addr_remain3_2668;
address_decode_4 decoder_3_2668 = address_decode_4(addr_selector2_166[12],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2668,addr_remain3_2668);


wire[15:0] addr_selector3_2669;
wire[15:0] addr_remain3_2669;
address_decode_4 decoder_3_2669 = address_decode_4(addr_selector2_166[13],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2669,addr_remain3_2669);


wire[15:0] addr_selector3_2670;
wire[15:0] addr_remain3_2670;
address_decode_4 decoder_3_2670 = address_decode_4(addr_selector2_166[14],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2670,addr_remain3_2670);


wire[15:0] addr_selector3_2671;
wire[15:0] addr_remain3_2671;
address_decode_4 decoder_3_2671 = address_decode_4(addr_selector2_166[15],addr_remain2_166[15:0],addr_remain2_166,addr_selector3_2671,addr_remain3_2671);


wire[15:0] addr_selector3_2672;
wire[15:0] addr_remain3_2672;
address_decode_4 decoder_3_2672 = address_decode_4(addr_selector2_167[0],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2672,addr_remain3_2672);


wire[15:0] addr_selector3_2673;
wire[15:0] addr_remain3_2673;
address_decode_4 decoder_3_2673 = address_decode_4(addr_selector2_167[1],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2673,addr_remain3_2673);


wire[15:0] addr_selector3_2674;
wire[15:0] addr_remain3_2674;
address_decode_4 decoder_3_2674 = address_decode_4(addr_selector2_167[2],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2674,addr_remain3_2674);


wire[15:0] addr_selector3_2675;
wire[15:0] addr_remain3_2675;
address_decode_4 decoder_3_2675 = address_decode_4(addr_selector2_167[3],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2675,addr_remain3_2675);


wire[15:0] addr_selector3_2676;
wire[15:0] addr_remain3_2676;
address_decode_4 decoder_3_2676 = address_decode_4(addr_selector2_167[4],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2676,addr_remain3_2676);


wire[15:0] addr_selector3_2677;
wire[15:0] addr_remain3_2677;
address_decode_4 decoder_3_2677 = address_decode_4(addr_selector2_167[5],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2677,addr_remain3_2677);


wire[15:0] addr_selector3_2678;
wire[15:0] addr_remain3_2678;
address_decode_4 decoder_3_2678 = address_decode_4(addr_selector2_167[6],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2678,addr_remain3_2678);


wire[15:0] addr_selector3_2679;
wire[15:0] addr_remain3_2679;
address_decode_4 decoder_3_2679 = address_decode_4(addr_selector2_167[7],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2679,addr_remain3_2679);


wire[15:0] addr_selector3_2680;
wire[15:0] addr_remain3_2680;
address_decode_4 decoder_3_2680 = address_decode_4(addr_selector2_167[8],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2680,addr_remain3_2680);


wire[15:0] addr_selector3_2681;
wire[15:0] addr_remain3_2681;
address_decode_4 decoder_3_2681 = address_decode_4(addr_selector2_167[9],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2681,addr_remain3_2681);


wire[15:0] addr_selector3_2682;
wire[15:0] addr_remain3_2682;
address_decode_4 decoder_3_2682 = address_decode_4(addr_selector2_167[10],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2682,addr_remain3_2682);


wire[15:0] addr_selector3_2683;
wire[15:0] addr_remain3_2683;
address_decode_4 decoder_3_2683 = address_decode_4(addr_selector2_167[11],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2683,addr_remain3_2683);


wire[15:0] addr_selector3_2684;
wire[15:0] addr_remain3_2684;
address_decode_4 decoder_3_2684 = address_decode_4(addr_selector2_167[12],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2684,addr_remain3_2684);


wire[15:0] addr_selector3_2685;
wire[15:0] addr_remain3_2685;
address_decode_4 decoder_3_2685 = address_decode_4(addr_selector2_167[13],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2685,addr_remain3_2685);


wire[15:0] addr_selector3_2686;
wire[15:0] addr_remain3_2686;
address_decode_4 decoder_3_2686 = address_decode_4(addr_selector2_167[14],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2686,addr_remain3_2686);


wire[15:0] addr_selector3_2687;
wire[15:0] addr_remain3_2687;
address_decode_4 decoder_3_2687 = address_decode_4(addr_selector2_167[15],addr_remain2_167[15:0],addr_remain2_167,addr_selector3_2687,addr_remain3_2687);


wire[15:0] addr_selector3_2688;
wire[15:0] addr_remain3_2688;
address_decode_4 decoder_3_2688 = address_decode_4(addr_selector2_168[0],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2688,addr_remain3_2688);


wire[15:0] addr_selector3_2689;
wire[15:0] addr_remain3_2689;
address_decode_4 decoder_3_2689 = address_decode_4(addr_selector2_168[1],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2689,addr_remain3_2689);


wire[15:0] addr_selector3_2690;
wire[15:0] addr_remain3_2690;
address_decode_4 decoder_3_2690 = address_decode_4(addr_selector2_168[2],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2690,addr_remain3_2690);


wire[15:0] addr_selector3_2691;
wire[15:0] addr_remain3_2691;
address_decode_4 decoder_3_2691 = address_decode_4(addr_selector2_168[3],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2691,addr_remain3_2691);


wire[15:0] addr_selector3_2692;
wire[15:0] addr_remain3_2692;
address_decode_4 decoder_3_2692 = address_decode_4(addr_selector2_168[4],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2692,addr_remain3_2692);


wire[15:0] addr_selector3_2693;
wire[15:0] addr_remain3_2693;
address_decode_4 decoder_3_2693 = address_decode_4(addr_selector2_168[5],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2693,addr_remain3_2693);


wire[15:0] addr_selector3_2694;
wire[15:0] addr_remain3_2694;
address_decode_4 decoder_3_2694 = address_decode_4(addr_selector2_168[6],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2694,addr_remain3_2694);


wire[15:0] addr_selector3_2695;
wire[15:0] addr_remain3_2695;
address_decode_4 decoder_3_2695 = address_decode_4(addr_selector2_168[7],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2695,addr_remain3_2695);


wire[15:0] addr_selector3_2696;
wire[15:0] addr_remain3_2696;
address_decode_4 decoder_3_2696 = address_decode_4(addr_selector2_168[8],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2696,addr_remain3_2696);


wire[15:0] addr_selector3_2697;
wire[15:0] addr_remain3_2697;
address_decode_4 decoder_3_2697 = address_decode_4(addr_selector2_168[9],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2697,addr_remain3_2697);


wire[15:0] addr_selector3_2698;
wire[15:0] addr_remain3_2698;
address_decode_4 decoder_3_2698 = address_decode_4(addr_selector2_168[10],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2698,addr_remain3_2698);


wire[15:0] addr_selector3_2699;
wire[15:0] addr_remain3_2699;
address_decode_4 decoder_3_2699 = address_decode_4(addr_selector2_168[11],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2699,addr_remain3_2699);


wire[15:0] addr_selector3_2700;
wire[15:0] addr_remain3_2700;
address_decode_4 decoder_3_2700 = address_decode_4(addr_selector2_168[12],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2700,addr_remain3_2700);


wire[15:0] addr_selector3_2701;
wire[15:0] addr_remain3_2701;
address_decode_4 decoder_3_2701 = address_decode_4(addr_selector2_168[13],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2701,addr_remain3_2701);


wire[15:0] addr_selector3_2702;
wire[15:0] addr_remain3_2702;
address_decode_4 decoder_3_2702 = address_decode_4(addr_selector2_168[14],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2702,addr_remain3_2702);


wire[15:0] addr_selector3_2703;
wire[15:0] addr_remain3_2703;
address_decode_4 decoder_3_2703 = address_decode_4(addr_selector2_168[15],addr_remain2_168[15:0],addr_remain2_168,addr_selector3_2703,addr_remain3_2703);


wire[15:0] addr_selector3_2704;
wire[15:0] addr_remain3_2704;
address_decode_4 decoder_3_2704 = address_decode_4(addr_selector2_169[0],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2704,addr_remain3_2704);


wire[15:0] addr_selector3_2705;
wire[15:0] addr_remain3_2705;
address_decode_4 decoder_3_2705 = address_decode_4(addr_selector2_169[1],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2705,addr_remain3_2705);


wire[15:0] addr_selector3_2706;
wire[15:0] addr_remain3_2706;
address_decode_4 decoder_3_2706 = address_decode_4(addr_selector2_169[2],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2706,addr_remain3_2706);


wire[15:0] addr_selector3_2707;
wire[15:0] addr_remain3_2707;
address_decode_4 decoder_3_2707 = address_decode_4(addr_selector2_169[3],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2707,addr_remain3_2707);


wire[15:0] addr_selector3_2708;
wire[15:0] addr_remain3_2708;
address_decode_4 decoder_3_2708 = address_decode_4(addr_selector2_169[4],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2708,addr_remain3_2708);


wire[15:0] addr_selector3_2709;
wire[15:0] addr_remain3_2709;
address_decode_4 decoder_3_2709 = address_decode_4(addr_selector2_169[5],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2709,addr_remain3_2709);


wire[15:0] addr_selector3_2710;
wire[15:0] addr_remain3_2710;
address_decode_4 decoder_3_2710 = address_decode_4(addr_selector2_169[6],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2710,addr_remain3_2710);


wire[15:0] addr_selector3_2711;
wire[15:0] addr_remain3_2711;
address_decode_4 decoder_3_2711 = address_decode_4(addr_selector2_169[7],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2711,addr_remain3_2711);


wire[15:0] addr_selector3_2712;
wire[15:0] addr_remain3_2712;
address_decode_4 decoder_3_2712 = address_decode_4(addr_selector2_169[8],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2712,addr_remain3_2712);


wire[15:0] addr_selector3_2713;
wire[15:0] addr_remain3_2713;
address_decode_4 decoder_3_2713 = address_decode_4(addr_selector2_169[9],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2713,addr_remain3_2713);


wire[15:0] addr_selector3_2714;
wire[15:0] addr_remain3_2714;
address_decode_4 decoder_3_2714 = address_decode_4(addr_selector2_169[10],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2714,addr_remain3_2714);


wire[15:0] addr_selector3_2715;
wire[15:0] addr_remain3_2715;
address_decode_4 decoder_3_2715 = address_decode_4(addr_selector2_169[11],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2715,addr_remain3_2715);


wire[15:0] addr_selector3_2716;
wire[15:0] addr_remain3_2716;
address_decode_4 decoder_3_2716 = address_decode_4(addr_selector2_169[12],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2716,addr_remain3_2716);


wire[15:0] addr_selector3_2717;
wire[15:0] addr_remain3_2717;
address_decode_4 decoder_3_2717 = address_decode_4(addr_selector2_169[13],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2717,addr_remain3_2717);


wire[15:0] addr_selector3_2718;
wire[15:0] addr_remain3_2718;
address_decode_4 decoder_3_2718 = address_decode_4(addr_selector2_169[14],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2718,addr_remain3_2718);


wire[15:0] addr_selector3_2719;
wire[15:0] addr_remain3_2719;
address_decode_4 decoder_3_2719 = address_decode_4(addr_selector2_169[15],addr_remain2_169[15:0],addr_remain2_169,addr_selector3_2719,addr_remain3_2719);


wire[15:0] addr_selector3_2720;
wire[15:0] addr_remain3_2720;
address_decode_4 decoder_3_2720 = address_decode_4(addr_selector2_170[0],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2720,addr_remain3_2720);


wire[15:0] addr_selector3_2721;
wire[15:0] addr_remain3_2721;
address_decode_4 decoder_3_2721 = address_decode_4(addr_selector2_170[1],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2721,addr_remain3_2721);


wire[15:0] addr_selector3_2722;
wire[15:0] addr_remain3_2722;
address_decode_4 decoder_3_2722 = address_decode_4(addr_selector2_170[2],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2722,addr_remain3_2722);


wire[15:0] addr_selector3_2723;
wire[15:0] addr_remain3_2723;
address_decode_4 decoder_3_2723 = address_decode_4(addr_selector2_170[3],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2723,addr_remain3_2723);


wire[15:0] addr_selector3_2724;
wire[15:0] addr_remain3_2724;
address_decode_4 decoder_3_2724 = address_decode_4(addr_selector2_170[4],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2724,addr_remain3_2724);


wire[15:0] addr_selector3_2725;
wire[15:0] addr_remain3_2725;
address_decode_4 decoder_3_2725 = address_decode_4(addr_selector2_170[5],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2725,addr_remain3_2725);


wire[15:0] addr_selector3_2726;
wire[15:0] addr_remain3_2726;
address_decode_4 decoder_3_2726 = address_decode_4(addr_selector2_170[6],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2726,addr_remain3_2726);


wire[15:0] addr_selector3_2727;
wire[15:0] addr_remain3_2727;
address_decode_4 decoder_3_2727 = address_decode_4(addr_selector2_170[7],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2727,addr_remain3_2727);


wire[15:0] addr_selector3_2728;
wire[15:0] addr_remain3_2728;
address_decode_4 decoder_3_2728 = address_decode_4(addr_selector2_170[8],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2728,addr_remain3_2728);


wire[15:0] addr_selector3_2729;
wire[15:0] addr_remain3_2729;
address_decode_4 decoder_3_2729 = address_decode_4(addr_selector2_170[9],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2729,addr_remain3_2729);


wire[15:0] addr_selector3_2730;
wire[15:0] addr_remain3_2730;
address_decode_4 decoder_3_2730 = address_decode_4(addr_selector2_170[10],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2730,addr_remain3_2730);


wire[15:0] addr_selector3_2731;
wire[15:0] addr_remain3_2731;
address_decode_4 decoder_3_2731 = address_decode_4(addr_selector2_170[11],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2731,addr_remain3_2731);


wire[15:0] addr_selector3_2732;
wire[15:0] addr_remain3_2732;
address_decode_4 decoder_3_2732 = address_decode_4(addr_selector2_170[12],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2732,addr_remain3_2732);


wire[15:0] addr_selector3_2733;
wire[15:0] addr_remain3_2733;
address_decode_4 decoder_3_2733 = address_decode_4(addr_selector2_170[13],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2733,addr_remain3_2733);


wire[15:0] addr_selector3_2734;
wire[15:0] addr_remain3_2734;
address_decode_4 decoder_3_2734 = address_decode_4(addr_selector2_170[14],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2734,addr_remain3_2734);


wire[15:0] addr_selector3_2735;
wire[15:0] addr_remain3_2735;
address_decode_4 decoder_3_2735 = address_decode_4(addr_selector2_170[15],addr_remain2_170[15:0],addr_remain2_170,addr_selector3_2735,addr_remain3_2735);


wire[15:0] addr_selector3_2736;
wire[15:0] addr_remain3_2736;
address_decode_4 decoder_3_2736 = address_decode_4(addr_selector2_171[0],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2736,addr_remain3_2736);


wire[15:0] addr_selector3_2737;
wire[15:0] addr_remain3_2737;
address_decode_4 decoder_3_2737 = address_decode_4(addr_selector2_171[1],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2737,addr_remain3_2737);


wire[15:0] addr_selector3_2738;
wire[15:0] addr_remain3_2738;
address_decode_4 decoder_3_2738 = address_decode_4(addr_selector2_171[2],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2738,addr_remain3_2738);


wire[15:0] addr_selector3_2739;
wire[15:0] addr_remain3_2739;
address_decode_4 decoder_3_2739 = address_decode_4(addr_selector2_171[3],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2739,addr_remain3_2739);


wire[15:0] addr_selector3_2740;
wire[15:0] addr_remain3_2740;
address_decode_4 decoder_3_2740 = address_decode_4(addr_selector2_171[4],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2740,addr_remain3_2740);


wire[15:0] addr_selector3_2741;
wire[15:0] addr_remain3_2741;
address_decode_4 decoder_3_2741 = address_decode_4(addr_selector2_171[5],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2741,addr_remain3_2741);


wire[15:0] addr_selector3_2742;
wire[15:0] addr_remain3_2742;
address_decode_4 decoder_3_2742 = address_decode_4(addr_selector2_171[6],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2742,addr_remain3_2742);


wire[15:0] addr_selector3_2743;
wire[15:0] addr_remain3_2743;
address_decode_4 decoder_3_2743 = address_decode_4(addr_selector2_171[7],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2743,addr_remain3_2743);


wire[15:0] addr_selector3_2744;
wire[15:0] addr_remain3_2744;
address_decode_4 decoder_3_2744 = address_decode_4(addr_selector2_171[8],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2744,addr_remain3_2744);


wire[15:0] addr_selector3_2745;
wire[15:0] addr_remain3_2745;
address_decode_4 decoder_3_2745 = address_decode_4(addr_selector2_171[9],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2745,addr_remain3_2745);


wire[15:0] addr_selector3_2746;
wire[15:0] addr_remain3_2746;
address_decode_4 decoder_3_2746 = address_decode_4(addr_selector2_171[10],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2746,addr_remain3_2746);


wire[15:0] addr_selector3_2747;
wire[15:0] addr_remain3_2747;
address_decode_4 decoder_3_2747 = address_decode_4(addr_selector2_171[11],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2747,addr_remain3_2747);


wire[15:0] addr_selector3_2748;
wire[15:0] addr_remain3_2748;
address_decode_4 decoder_3_2748 = address_decode_4(addr_selector2_171[12],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2748,addr_remain3_2748);


wire[15:0] addr_selector3_2749;
wire[15:0] addr_remain3_2749;
address_decode_4 decoder_3_2749 = address_decode_4(addr_selector2_171[13],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2749,addr_remain3_2749);


wire[15:0] addr_selector3_2750;
wire[15:0] addr_remain3_2750;
address_decode_4 decoder_3_2750 = address_decode_4(addr_selector2_171[14],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2750,addr_remain3_2750);


wire[15:0] addr_selector3_2751;
wire[15:0] addr_remain3_2751;
address_decode_4 decoder_3_2751 = address_decode_4(addr_selector2_171[15],addr_remain2_171[15:0],addr_remain2_171,addr_selector3_2751,addr_remain3_2751);


wire[15:0] addr_selector3_2752;
wire[15:0] addr_remain3_2752;
address_decode_4 decoder_3_2752 = address_decode_4(addr_selector2_172[0],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2752,addr_remain3_2752);


wire[15:0] addr_selector3_2753;
wire[15:0] addr_remain3_2753;
address_decode_4 decoder_3_2753 = address_decode_4(addr_selector2_172[1],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2753,addr_remain3_2753);


wire[15:0] addr_selector3_2754;
wire[15:0] addr_remain3_2754;
address_decode_4 decoder_3_2754 = address_decode_4(addr_selector2_172[2],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2754,addr_remain3_2754);


wire[15:0] addr_selector3_2755;
wire[15:0] addr_remain3_2755;
address_decode_4 decoder_3_2755 = address_decode_4(addr_selector2_172[3],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2755,addr_remain3_2755);


wire[15:0] addr_selector3_2756;
wire[15:0] addr_remain3_2756;
address_decode_4 decoder_3_2756 = address_decode_4(addr_selector2_172[4],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2756,addr_remain3_2756);


wire[15:0] addr_selector3_2757;
wire[15:0] addr_remain3_2757;
address_decode_4 decoder_3_2757 = address_decode_4(addr_selector2_172[5],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2757,addr_remain3_2757);


wire[15:0] addr_selector3_2758;
wire[15:0] addr_remain3_2758;
address_decode_4 decoder_3_2758 = address_decode_4(addr_selector2_172[6],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2758,addr_remain3_2758);


wire[15:0] addr_selector3_2759;
wire[15:0] addr_remain3_2759;
address_decode_4 decoder_3_2759 = address_decode_4(addr_selector2_172[7],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2759,addr_remain3_2759);


wire[15:0] addr_selector3_2760;
wire[15:0] addr_remain3_2760;
address_decode_4 decoder_3_2760 = address_decode_4(addr_selector2_172[8],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2760,addr_remain3_2760);


wire[15:0] addr_selector3_2761;
wire[15:0] addr_remain3_2761;
address_decode_4 decoder_3_2761 = address_decode_4(addr_selector2_172[9],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2761,addr_remain3_2761);


wire[15:0] addr_selector3_2762;
wire[15:0] addr_remain3_2762;
address_decode_4 decoder_3_2762 = address_decode_4(addr_selector2_172[10],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2762,addr_remain3_2762);


wire[15:0] addr_selector3_2763;
wire[15:0] addr_remain3_2763;
address_decode_4 decoder_3_2763 = address_decode_4(addr_selector2_172[11],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2763,addr_remain3_2763);


wire[15:0] addr_selector3_2764;
wire[15:0] addr_remain3_2764;
address_decode_4 decoder_3_2764 = address_decode_4(addr_selector2_172[12],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2764,addr_remain3_2764);


wire[15:0] addr_selector3_2765;
wire[15:0] addr_remain3_2765;
address_decode_4 decoder_3_2765 = address_decode_4(addr_selector2_172[13],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2765,addr_remain3_2765);


wire[15:0] addr_selector3_2766;
wire[15:0] addr_remain3_2766;
address_decode_4 decoder_3_2766 = address_decode_4(addr_selector2_172[14],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2766,addr_remain3_2766);


wire[15:0] addr_selector3_2767;
wire[15:0] addr_remain3_2767;
address_decode_4 decoder_3_2767 = address_decode_4(addr_selector2_172[15],addr_remain2_172[15:0],addr_remain2_172,addr_selector3_2767,addr_remain3_2767);


wire[15:0] addr_selector3_2768;
wire[15:0] addr_remain3_2768;
address_decode_4 decoder_3_2768 = address_decode_4(addr_selector2_173[0],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2768,addr_remain3_2768);


wire[15:0] addr_selector3_2769;
wire[15:0] addr_remain3_2769;
address_decode_4 decoder_3_2769 = address_decode_4(addr_selector2_173[1],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2769,addr_remain3_2769);


wire[15:0] addr_selector3_2770;
wire[15:0] addr_remain3_2770;
address_decode_4 decoder_3_2770 = address_decode_4(addr_selector2_173[2],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2770,addr_remain3_2770);


wire[15:0] addr_selector3_2771;
wire[15:0] addr_remain3_2771;
address_decode_4 decoder_3_2771 = address_decode_4(addr_selector2_173[3],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2771,addr_remain3_2771);


wire[15:0] addr_selector3_2772;
wire[15:0] addr_remain3_2772;
address_decode_4 decoder_3_2772 = address_decode_4(addr_selector2_173[4],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2772,addr_remain3_2772);


wire[15:0] addr_selector3_2773;
wire[15:0] addr_remain3_2773;
address_decode_4 decoder_3_2773 = address_decode_4(addr_selector2_173[5],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2773,addr_remain3_2773);


wire[15:0] addr_selector3_2774;
wire[15:0] addr_remain3_2774;
address_decode_4 decoder_3_2774 = address_decode_4(addr_selector2_173[6],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2774,addr_remain3_2774);


wire[15:0] addr_selector3_2775;
wire[15:0] addr_remain3_2775;
address_decode_4 decoder_3_2775 = address_decode_4(addr_selector2_173[7],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2775,addr_remain3_2775);


wire[15:0] addr_selector3_2776;
wire[15:0] addr_remain3_2776;
address_decode_4 decoder_3_2776 = address_decode_4(addr_selector2_173[8],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2776,addr_remain3_2776);


wire[15:0] addr_selector3_2777;
wire[15:0] addr_remain3_2777;
address_decode_4 decoder_3_2777 = address_decode_4(addr_selector2_173[9],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2777,addr_remain3_2777);


wire[15:0] addr_selector3_2778;
wire[15:0] addr_remain3_2778;
address_decode_4 decoder_3_2778 = address_decode_4(addr_selector2_173[10],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2778,addr_remain3_2778);


wire[15:0] addr_selector3_2779;
wire[15:0] addr_remain3_2779;
address_decode_4 decoder_3_2779 = address_decode_4(addr_selector2_173[11],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2779,addr_remain3_2779);


wire[15:0] addr_selector3_2780;
wire[15:0] addr_remain3_2780;
address_decode_4 decoder_3_2780 = address_decode_4(addr_selector2_173[12],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2780,addr_remain3_2780);


wire[15:0] addr_selector3_2781;
wire[15:0] addr_remain3_2781;
address_decode_4 decoder_3_2781 = address_decode_4(addr_selector2_173[13],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2781,addr_remain3_2781);


wire[15:0] addr_selector3_2782;
wire[15:0] addr_remain3_2782;
address_decode_4 decoder_3_2782 = address_decode_4(addr_selector2_173[14],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2782,addr_remain3_2782);


wire[15:0] addr_selector3_2783;
wire[15:0] addr_remain3_2783;
address_decode_4 decoder_3_2783 = address_decode_4(addr_selector2_173[15],addr_remain2_173[15:0],addr_remain2_173,addr_selector3_2783,addr_remain3_2783);


wire[15:0] addr_selector3_2784;
wire[15:0] addr_remain3_2784;
address_decode_4 decoder_3_2784 = address_decode_4(addr_selector2_174[0],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2784,addr_remain3_2784);


wire[15:0] addr_selector3_2785;
wire[15:0] addr_remain3_2785;
address_decode_4 decoder_3_2785 = address_decode_4(addr_selector2_174[1],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2785,addr_remain3_2785);


wire[15:0] addr_selector3_2786;
wire[15:0] addr_remain3_2786;
address_decode_4 decoder_3_2786 = address_decode_4(addr_selector2_174[2],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2786,addr_remain3_2786);


wire[15:0] addr_selector3_2787;
wire[15:0] addr_remain3_2787;
address_decode_4 decoder_3_2787 = address_decode_4(addr_selector2_174[3],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2787,addr_remain3_2787);


wire[15:0] addr_selector3_2788;
wire[15:0] addr_remain3_2788;
address_decode_4 decoder_3_2788 = address_decode_4(addr_selector2_174[4],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2788,addr_remain3_2788);


wire[15:0] addr_selector3_2789;
wire[15:0] addr_remain3_2789;
address_decode_4 decoder_3_2789 = address_decode_4(addr_selector2_174[5],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2789,addr_remain3_2789);


wire[15:0] addr_selector3_2790;
wire[15:0] addr_remain3_2790;
address_decode_4 decoder_3_2790 = address_decode_4(addr_selector2_174[6],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2790,addr_remain3_2790);


wire[15:0] addr_selector3_2791;
wire[15:0] addr_remain3_2791;
address_decode_4 decoder_3_2791 = address_decode_4(addr_selector2_174[7],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2791,addr_remain3_2791);


wire[15:0] addr_selector3_2792;
wire[15:0] addr_remain3_2792;
address_decode_4 decoder_3_2792 = address_decode_4(addr_selector2_174[8],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2792,addr_remain3_2792);


wire[15:0] addr_selector3_2793;
wire[15:0] addr_remain3_2793;
address_decode_4 decoder_3_2793 = address_decode_4(addr_selector2_174[9],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2793,addr_remain3_2793);


wire[15:0] addr_selector3_2794;
wire[15:0] addr_remain3_2794;
address_decode_4 decoder_3_2794 = address_decode_4(addr_selector2_174[10],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2794,addr_remain3_2794);


wire[15:0] addr_selector3_2795;
wire[15:0] addr_remain3_2795;
address_decode_4 decoder_3_2795 = address_decode_4(addr_selector2_174[11],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2795,addr_remain3_2795);


wire[15:0] addr_selector3_2796;
wire[15:0] addr_remain3_2796;
address_decode_4 decoder_3_2796 = address_decode_4(addr_selector2_174[12],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2796,addr_remain3_2796);


wire[15:0] addr_selector3_2797;
wire[15:0] addr_remain3_2797;
address_decode_4 decoder_3_2797 = address_decode_4(addr_selector2_174[13],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2797,addr_remain3_2797);


wire[15:0] addr_selector3_2798;
wire[15:0] addr_remain3_2798;
address_decode_4 decoder_3_2798 = address_decode_4(addr_selector2_174[14],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2798,addr_remain3_2798);


wire[15:0] addr_selector3_2799;
wire[15:0] addr_remain3_2799;
address_decode_4 decoder_3_2799 = address_decode_4(addr_selector2_174[15],addr_remain2_174[15:0],addr_remain2_174,addr_selector3_2799,addr_remain3_2799);


wire[15:0] addr_selector3_2800;
wire[15:0] addr_remain3_2800;
address_decode_4 decoder_3_2800 = address_decode_4(addr_selector2_175[0],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2800,addr_remain3_2800);


wire[15:0] addr_selector3_2801;
wire[15:0] addr_remain3_2801;
address_decode_4 decoder_3_2801 = address_decode_4(addr_selector2_175[1],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2801,addr_remain3_2801);


wire[15:0] addr_selector3_2802;
wire[15:0] addr_remain3_2802;
address_decode_4 decoder_3_2802 = address_decode_4(addr_selector2_175[2],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2802,addr_remain3_2802);


wire[15:0] addr_selector3_2803;
wire[15:0] addr_remain3_2803;
address_decode_4 decoder_3_2803 = address_decode_4(addr_selector2_175[3],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2803,addr_remain3_2803);


wire[15:0] addr_selector3_2804;
wire[15:0] addr_remain3_2804;
address_decode_4 decoder_3_2804 = address_decode_4(addr_selector2_175[4],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2804,addr_remain3_2804);


wire[15:0] addr_selector3_2805;
wire[15:0] addr_remain3_2805;
address_decode_4 decoder_3_2805 = address_decode_4(addr_selector2_175[5],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2805,addr_remain3_2805);


wire[15:0] addr_selector3_2806;
wire[15:0] addr_remain3_2806;
address_decode_4 decoder_3_2806 = address_decode_4(addr_selector2_175[6],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2806,addr_remain3_2806);


wire[15:0] addr_selector3_2807;
wire[15:0] addr_remain3_2807;
address_decode_4 decoder_3_2807 = address_decode_4(addr_selector2_175[7],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2807,addr_remain3_2807);


wire[15:0] addr_selector3_2808;
wire[15:0] addr_remain3_2808;
address_decode_4 decoder_3_2808 = address_decode_4(addr_selector2_175[8],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2808,addr_remain3_2808);


wire[15:0] addr_selector3_2809;
wire[15:0] addr_remain3_2809;
address_decode_4 decoder_3_2809 = address_decode_4(addr_selector2_175[9],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2809,addr_remain3_2809);


wire[15:0] addr_selector3_2810;
wire[15:0] addr_remain3_2810;
address_decode_4 decoder_3_2810 = address_decode_4(addr_selector2_175[10],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2810,addr_remain3_2810);


wire[15:0] addr_selector3_2811;
wire[15:0] addr_remain3_2811;
address_decode_4 decoder_3_2811 = address_decode_4(addr_selector2_175[11],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2811,addr_remain3_2811);


wire[15:0] addr_selector3_2812;
wire[15:0] addr_remain3_2812;
address_decode_4 decoder_3_2812 = address_decode_4(addr_selector2_175[12],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2812,addr_remain3_2812);


wire[15:0] addr_selector3_2813;
wire[15:0] addr_remain3_2813;
address_decode_4 decoder_3_2813 = address_decode_4(addr_selector2_175[13],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2813,addr_remain3_2813);


wire[15:0] addr_selector3_2814;
wire[15:0] addr_remain3_2814;
address_decode_4 decoder_3_2814 = address_decode_4(addr_selector2_175[14],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2814,addr_remain3_2814);


wire[15:0] addr_selector3_2815;
wire[15:0] addr_remain3_2815;
address_decode_4 decoder_3_2815 = address_decode_4(addr_selector2_175[15],addr_remain2_175[15:0],addr_remain2_175,addr_selector3_2815,addr_remain3_2815);


wire[15:0] addr_selector3_2816;
wire[15:0] addr_remain3_2816;
address_decode_4 decoder_3_2816 = address_decode_4(addr_selector2_176[0],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2816,addr_remain3_2816);


wire[15:0] addr_selector3_2817;
wire[15:0] addr_remain3_2817;
address_decode_4 decoder_3_2817 = address_decode_4(addr_selector2_176[1],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2817,addr_remain3_2817);


wire[15:0] addr_selector3_2818;
wire[15:0] addr_remain3_2818;
address_decode_4 decoder_3_2818 = address_decode_4(addr_selector2_176[2],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2818,addr_remain3_2818);


wire[15:0] addr_selector3_2819;
wire[15:0] addr_remain3_2819;
address_decode_4 decoder_3_2819 = address_decode_4(addr_selector2_176[3],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2819,addr_remain3_2819);


wire[15:0] addr_selector3_2820;
wire[15:0] addr_remain3_2820;
address_decode_4 decoder_3_2820 = address_decode_4(addr_selector2_176[4],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2820,addr_remain3_2820);


wire[15:0] addr_selector3_2821;
wire[15:0] addr_remain3_2821;
address_decode_4 decoder_3_2821 = address_decode_4(addr_selector2_176[5],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2821,addr_remain3_2821);


wire[15:0] addr_selector3_2822;
wire[15:0] addr_remain3_2822;
address_decode_4 decoder_3_2822 = address_decode_4(addr_selector2_176[6],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2822,addr_remain3_2822);


wire[15:0] addr_selector3_2823;
wire[15:0] addr_remain3_2823;
address_decode_4 decoder_3_2823 = address_decode_4(addr_selector2_176[7],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2823,addr_remain3_2823);


wire[15:0] addr_selector3_2824;
wire[15:0] addr_remain3_2824;
address_decode_4 decoder_3_2824 = address_decode_4(addr_selector2_176[8],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2824,addr_remain3_2824);


wire[15:0] addr_selector3_2825;
wire[15:0] addr_remain3_2825;
address_decode_4 decoder_3_2825 = address_decode_4(addr_selector2_176[9],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2825,addr_remain3_2825);


wire[15:0] addr_selector3_2826;
wire[15:0] addr_remain3_2826;
address_decode_4 decoder_3_2826 = address_decode_4(addr_selector2_176[10],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2826,addr_remain3_2826);


wire[15:0] addr_selector3_2827;
wire[15:0] addr_remain3_2827;
address_decode_4 decoder_3_2827 = address_decode_4(addr_selector2_176[11],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2827,addr_remain3_2827);


wire[15:0] addr_selector3_2828;
wire[15:0] addr_remain3_2828;
address_decode_4 decoder_3_2828 = address_decode_4(addr_selector2_176[12],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2828,addr_remain3_2828);


wire[15:0] addr_selector3_2829;
wire[15:0] addr_remain3_2829;
address_decode_4 decoder_3_2829 = address_decode_4(addr_selector2_176[13],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2829,addr_remain3_2829);


wire[15:0] addr_selector3_2830;
wire[15:0] addr_remain3_2830;
address_decode_4 decoder_3_2830 = address_decode_4(addr_selector2_176[14],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2830,addr_remain3_2830);


wire[15:0] addr_selector3_2831;
wire[15:0] addr_remain3_2831;
address_decode_4 decoder_3_2831 = address_decode_4(addr_selector2_176[15],addr_remain2_176[15:0],addr_remain2_176,addr_selector3_2831,addr_remain3_2831);


wire[15:0] addr_selector3_2832;
wire[15:0] addr_remain3_2832;
address_decode_4 decoder_3_2832 = address_decode_4(addr_selector2_177[0],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2832,addr_remain3_2832);


wire[15:0] addr_selector3_2833;
wire[15:0] addr_remain3_2833;
address_decode_4 decoder_3_2833 = address_decode_4(addr_selector2_177[1],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2833,addr_remain3_2833);


wire[15:0] addr_selector3_2834;
wire[15:0] addr_remain3_2834;
address_decode_4 decoder_3_2834 = address_decode_4(addr_selector2_177[2],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2834,addr_remain3_2834);


wire[15:0] addr_selector3_2835;
wire[15:0] addr_remain3_2835;
address_decode_4 decoder_3_2835 = address_decode_4(addr_selector2_177[3],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2835,addr_remain3_2835);


wire[15:0] addr_selector3_2836;
wire[15:0] addr_remain3_2836;
address_decode_4 decoder_3_2836 = address_decode_4(addr_selector2_177[4],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2836,addr_remain3_2836);


wire[15:0] addr_selector3_2837;
wire[15:0] addr_remain3_2837;
address_decode_4 decoder_3_2837 = address_decode_4(addr_selector2_177[5],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2837,addr_remain3_2837);


wire[15:0] addr_selector3_2838;
wire[15:0] addr_remain3_2838;
address_decode_4 decoder_3_2838 = address_decode_4(addr_selector2_177[6],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2838,addr_remain3_2838);


wire[15:0] addr_selector3_2839;
wire[15:0] addr_remain3_2839;
address_decode_4 decoder_3_2839 = address_decode_4(addr_selector2_177[7],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2839,addr_remain3_2839);


wire[15:0] addr_selector3_2840;
wire[15:0] addr_remain3_2840;
address_decode_4 decoder_3_2840 = address_decode_4(addr_selector2_177[8],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2840,addr_remain3_2840);


wire[15:0] addr_selector3_2841;
wire[15:0] addr_remain3_2841;
address_decode_4 decoder_3_2841 = address_decode_4(addr_selector2_177[9],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2841,addr_remain3_2841);


wire[15:0] addr_selector3_2842;
wire[15:0] addr_remain3_2842;
address_decode_4 decoder_3_2842 = address_decode_4(addr_selector2_177[10],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2842,addr_remain3_2842);


wire[15:0] addr_selector3_2843;
wire[15:0] addr_remain3_2843;
address_decode_4 decoder_3_2843 = address_decode_4(addr_selector2_177[11],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2843,addr_remain3_2843);


wire[15:0] addr_selector3_2844;
wire[15:0] addr_remain3_2844;
address_decode_4 decoder_3_2844 = address_decode_4(addr_selector2_177[12],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2844,addr_remain3_2844);


wire[15:0] addr_selector3_2845;
wire[15:0] addr_remain3_2845;
address_decode_4 decoder_3_2845 = address_decode_4(addr_selector2_177[13],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2845,addr_remain3_2845);


wire[15:0] addr_selector3_2846;
wire[15:0] addr_remain3_2846;
address_decode_4 decoder_3_2846 = address_decode_4(addr_selector2_177[14],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2846,addr_remain3_2846);


wire[15:0] addr_selector3_2847;
wire[15:0] addr_remain3_2847;
address_decode_4 decoder_3_2847 = address_decode_4(addr_selector2_177[15],addr_remain2_177[15:0],addr_remain2_177,addr_selector3_2847,addr_remain3_2847);


wire[15:0] addr_selector3_2848;
wire[15:0] addr_remain3_2848;
address_decode_4 decoder_3_2848 = address_decode_4(addr_selector2_178[0],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2848,addr_remain3_2848);


wire[15:0] addr_selector3_2849;
wire[15:0] addr_remain3_2849;
address_decode_4 decoder_3_2849 = address_decode_4(addr_selector2_178[1],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2849,addr_remain3_2849);


wire[15:0] addr_selector3_2850;
wire[15:0] addr_remain3_2850;
address_decode_4 decoder_3_2850 = address_decode_4(addr_selector2_178[2],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2850,addr_remain3_2850);


wire[15:0] addr_selector3_2851;
wire[15:0] addr_remain3_2851;
address_decode_4 decoder_3_2851 = address_decode_4(addr_selector2_178[3],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2851,addr_remain3_2851);


wire[15:0] addr_selector3_2852;
wire[15:0] addr_remain3_2852;
address_decode_4 decoder_3_2852 = address_decode_4(addr_selector2_178[4],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2852,addr_remain3_2852);


wire[15:0] addr_selector3_2853;
wire[15:0] addr_remain3_2853;
address_decode_4 decoder_3_2853 = address_decode_4(addr_selector2_178[5],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2853,addr_remain3_2853);


wire[15:0] addr_selector3_2854;
wire[15:0] addr_remain3_2854;
address_decode_4 decoder_3_2854 = address_decode_4(addr_selector2_178[6],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2854,addr_remain3_2854);


wire[15:0] addr_selector3_2855;
wire[15:0] addr_remain3_2855;
address_decode_4 decoder_3_2855 = address_decode_4(addr_selector2_178[7],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2855,addr_remain3_2855);


wire[15:0] addr_selector3_2856;
wire[15:0] addr_remain3_2856;
address_decode_4 decoder_3_2856 = address_decode_4(addr_selector2_178[8],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2856,addr_remain3_2856);


wire[15:0] addr_selector3_2857;
wire[15:0] addr_remain3_2857;
address_decode_4 decoder_3_2857 = address_decode_4(addr_selector2_178[9],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2857,addr_remain3_2857);


wire[15:0] addr_selector3_2858;
wire[15:0] addr_remain3_2858;
address_decode_4 decoder_3_2858 = address_decode_4(addr_selector2_178[10],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2858,addr_remain3_2858);


wire[15:0] addr_selector3_2859;
wire[15:0] addr_remain3_2859;
address_decode_4 decoder_3_2859 = address_decode_4(addr_selector2_178[11],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2859,addr_remain3_2859);


wire[15:0] addr_selector3_2860;
wire[15:0] addr_remain3_2860;
address_decode_4 decoder_3_2860 = address_decode_4(addr_selector2_178[12],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2860,addr_remain3_2860);


wire[15:0] addr_selector3_2861;
wire[15:0] addr_remain3_2861;
address_decode_4 decoder_3_2861 = address_decode_4(addr_selector2_178[13],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2861,addr_remain3_2861);


wire[15:0] addr_selector3_2862;
wire[15:0] addr_remain3_2862;
address_decode_4 decoder_3_2862 = address_decode_4(addr_selector2_178[14],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2862,addr_remain3_2862);


wire[15:0] addr_selector3_2863;
wire[15:0] addr_remain3_2863;
address_decode_4 decoder_3_2863 = address_decode_4(addr_selector2_178[15],addr_remain2_178[15:0],addr_remain2_178,addr_selector3_2863,addr_remain3_2863);


wire[15:0] addr_selector3_2864;
wire[15:0] addr_remain3_2864;
address_decode_4 decoder_3_2864 = address_decode_4(addr_selector2_179[0],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2864,addr_remain3_2864);


wire[15:0] addr_selector3_2865;
wire[15:0] addr_remain3_2865;
address_decode_4 decoder_3_2865 = address_decode_4(addr_selector2_179[1],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2865,addr_remain3_2865);


wire[15:0] addr_selector3_2866;
wire[15:0] addr_remain3_2866;
address_decode_4 decoder_3_2866 = address_decode_4(addr_selector2_179[2],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2866,addr_remain3_2866);


wire[15:0] addr_selector3_2867;
wire[15:0] addr_remain3_2867;
address_decode_4 decoder_3_2867 = address_decode_4(addr_selector2_179[3],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2867,addr_remain3_2867);


wire[15:0] addr_selector3_2868;
wire[15:0] addr_remain3_2868;
address_decode_4 decoder_3_2868 = address_decode_4(addr_selector2_179[4],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2868,addr_remain3_2868);


wire[15:0] addr_selector3_2869;
wire[15:0] addr_remain3_2869;
address_decode_4 decoder_3_2869 = address_decode_4(addr_selector2_179[5],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2869,addr_remain3_2869);


wire[15:0] addr_selector3_2870;
wire[15:0] addr_remain3_2870;
address_decode_4 decoder_3_2870 = address_decode_4(addr_selector2_179[6],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2870,addr_remain3_2870);


wire[15:0] addr_selector3_2871;
wire[15:0] addr_remain3_2871;
address_decode_4 decoder_3_2871 = address_decode_4(addr_selector2_179[7],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2871,addr_remain3_2871);


wire[15:0] addr_selector3_2872;
wire[15:0] addr_remain3_2872;
address_decode_4 decoder_3_2872 = address_decode_4(addr_selector2_179[8],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2872,addr_remain3_2872);


wire[15:0] addr_selector3_2873;
wire[15:0] addr_remain3_2873;
address_decode_4 decoder_3_2873 = address_decode_4(addr_selector2_179[9],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2873,addr_remain3_2873);


wire[15:0] addr_selector3_2874;
wire[15:0] addr_remain3_2874;
address_decode_4 decoder_3_2874 = address_decode_4(addr_selector2_179[10],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2874,addr_remain3_2874);


wire[15:0] addr_selector3_2875;
wire[15:0] addr_remain3_2875;
address_decode_4 decoder_3_2875 = address_decode_4(addr_selector2_179[11],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2875,addr_remain3_2875);


wire[15:0] addr_selector3_2876;
wire[15:0] addr_remain3_2876;
address_decode_4 decoder_3_2876 = address_decode_4(addr_selector2_179[12],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2876,addr_remain3_2876);


wire[15:0] addr_selector3_2877;
wire[15:0] addr_remain3_2877;
address_decode_4 decoder_3_2877 = address_decode_4(addr_selector2_179[13],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2877,addr_remain3_2877);


wire[15:0] addr_selector3_2878;
wire[15:0] addr_remain3_2878;
address_decode_4 decoder_3_2878 = address_decode_4(addr_selector2_179[14],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2878,addr_remain3_2878);


wire[15:0] addr_selector3_2879;
wire[15:0] addr_remain3_2879;
address_decode_4 decoder_3_2879 = address_decode_4(addr_selector2_179[15],addr_remain2_179[15:0],addr_remain2_179,addr_selector3_2879,addr_remain3_2879);


wire[15:0] addr_selector3_2880;
wire[15:0] addr_remain3_2880;
address_decode_4 decoder_3_2880 = address_decode_4(addr_selector2_180[0],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2880,addr_remain3_2880);


wire[15:0] addr_selector3_2881;
wire[15:0] addr_remain3_2881;
address_decode_4 decoder_3_2881 = address_decode_4(addr_selector2_180[1],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2881,addr_remain3_2881);


wire[15:0] addr_selector3_2882;
wire[15:0] addr_remain3_2882;
address_decode_4 decoder_3_2882 = address_decode_4(addr_selector2_180[2],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2882,addr_remain3_2882);


wire[15:0] addr_selector3_2883;
wire[15:0] addr_remain3_2883;
address_decode_4 decoder_3_2883 = address_decode_4(addr_selector2_180[3],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2883,addr_remain3_2883);


wire[15:0] addr_selector3_2884;
wire[15:0] addr_remain3_2884;
address_decode_4 decoder_3_2884 = address_decode_4(addr_selector2_180[4],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2884,addr_remain3_2884);


wire[15:0] addr_selector3_2885;
wire[15:0] addr_remain3_2885;
address_decode_4 decoder_3_2885 = address_decode_4(addr_selector2_180[5],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2885,addr_remain3_2885);


wire[15:0] addr_selector3_2886;
wire[15:0] addr_remain3_2886;
address_decode_4 decoder_3_2886 = address_decode_4(addr_selector2_180[6],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2886,addr_remain3_2886);


wire[15:0] addr_selector3_2887;
wire[15:0] addr_remain3_2887;
address_decode_4 decoder_3_2887 = address_decode_4(addr_selector2_180[7],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2887,addr_remain3_2887);


wire[15:0] addr_selector3_2888;
wire[15:0] addr_remain3_2888;
address_decode_4 decoder_3_2888 = address_decode_4(addr_selector2_180[8],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2888,addr_remain3_2888);


wire[15:0] addr_selector3_2889;
wire[15:0] addr_remain3_2889;
address_decode_4 decoder_3_2889 = address_decode_4(addr_selector2_180[9],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2889,addr_remain3_2889);


wire[15:0] addr_selector3_2890;
wire[15:0] addr_remain3_2890;
address_decode_4 decoder_3_2890 = address_decode_4(addr_selector2_180[10],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2890,addr_remain3_2890);


wire[15:0] addr_selector3_2891;
wire[15:0] addr_remain3_2891;
address_decode_4 decoder_3_2891 = address_decode_4(addr_selector2_180[11],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2891,addr_remain3_2891);


wire[15:0] addr_selector3_2892;
wire[15:0] addr_remain3_2892;
address_decode_4 decoder_3_2892 = address_decode_4(addr_selector2_180[12],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2892,addr_remain3_2892);


wire[15:0] addr_selector3_2893;
wire[15:0] addr_remain3_2893;
address_decode_4 decoder_3_2893 = address_decode_4(addr_selector2_180[13],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2893,addr_remain3_2893);


wire[15:0] addr_selector3_2894;
wire[15:0] addr_remain3_2894;
address_decode_4 decoder_3_2894 = address_decode_4(addr_selector2_180[14],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2894,addr_remain3_2894);


wire[15:0] addr_selector3_2895;
wire[15:0] addr_remain3_2895;
address_decode_4 decoder_3_2895 = address_decode_4(addr_selector2_180[15],addr_remain2_180[15:0],addr_remain2_180,addr_selector3_2895,addr_remain3_2895);


wire[15:0] addr_selector3_2896;
wire[15:0] addr_remain3_2896;
address_decode_4 decoder_3_2896 = address_decode_4(addr_selector2_181[0],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2896,addr_remain3_2896);


wire[15:0] addr_selector3_2897;
wire[15:0] addr_remain3_2897;
address_decode_4 decoder_3_2897 = address_decode_4(addr_selector2_181[1],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2897,addr_remain3_2897);


wire[15:0] addr_selector3_2898;
wire[15:0] addr_remain3_2898;
address_decode_4 decoder_3_2898 = address_decode_4(addr_selector2_181[2],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2898,addr_remain3_2898);


wire[15:0] addr_selector3_2899;
wire[15:0] addr_remain3_2899;
address_decode_4 decoder_3_2899 = address_decode_4(addr_selector2_181[3],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2899,addr_remain3_2899);


wire[15:0] addr_selector3_2900;
wire[15:0] addr_remain3_2900;
address_decode_4 decoder_3_2900 = address_decode_4(addr_selector2_181[4],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2900,addr_remain3_2900);


wire[15:0] addr_selector3_2901;
wire[15:0] addr_remain3_2901;
address_decode_4 decoder_3_2901 = address_decode_4(addr_selector2_181[5],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2901,addr_remain3_2901);


wire[15:0] addr_selector3_2902;
wire[15:0] addr_remain3_2902;
address_decode_4 decoder_3_2902 = address_decode_4(addr_selector2_181[6],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2902,addr_remain3_2902);


wire[15:0] addr_selector3_2903;
wire[15:0] addr_remain3_2903;
address_decode_4 decoder_3_2903 = address_decode_4(addr_selector2_181[7],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2903,addr_remain3_2903);


wire[15:0] addr_selector3_2904;
wire[15:0] addr_remain3_2904;
address_decode_4 decoder_3_2904 = address_decode_4(addr_selector2_181[8],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2904,addr_remain3_2904);


wire[15:0] addr_selector3_2905;
wire[15:0] addr_remain3_2905;
address_decode_4 decoder_3_2905 = address_decode_4(addr_selector2_181[9],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2905,addr_remain3_2905);


wire[15:0] addr_selector3_2906;
wire[15:0] addr_remain3_2906;
address_decode_4 decoder_3_2906 = address_decode_4(addr_selector2_181[10],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2906,addr_remain3_2906);


wire[15:0] addr_selector3_2907;
wire[15:0] addr_remain3_2907;
address_decode_4 decoder_3_2907 = address_decode_4(addr_selector2_181[11],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2907,addr_remain3_2907);


wire[15:0] addr_selector3_2908;
wire[15:0] addr_remain3_2908;
address_decode_4 decoder_3_2908 = address_decode_4(addr_selector2_181[12],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2908,addr_remain3_2908);


wire[15:0] addr_selector3_2909;
wire[15:0] addr_remain3_2909;
address_decode_4 decoder_3_2909 = address_decode_4(addr_selector2_181[13],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2909,addr_remain3_2909);


wire[15:0] addr_selector3_2910;
wire[15:0] addr_remain3_2910;
address_decode_4 decoder_3_2910 = address_decode_4(addr_selector2_181[14],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2910,addr_remain3_2910);


wire[15:0] addr_selector3_2911;
wire[15:0] addr_remain3_2911;
address_decode_4 decoder_3_2911 = address_decode_4(addr_selector2_181[15],addr_remain2_181[15:0],addr_remain2_181,addr_selector3_2911,addr_remain3_2911);


wire[15:0] addr_selector3_2912;
wire[15:0] addr_remain3_2912;
address_decode_4 decoder_3_2912 = address_decode_4(addr_selector2_182[0],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2912,addr_remain3_2912);


wire[15:0] addr_selector3_2913;
wire[15:0] addr_remain3_2913;
address_decode_4 decoder_3_2913 = address_decode_4(addr_selector2_182[1],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2913,addr_remain3_2913);


wire[15:0] addr_selector3_2914;
wire[15:0] addr_remain3_2914;
address_decode_4 decoder_3_2914 = address_decode_4(addr_selector2_182[2],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2914,addr_remain3_2914);


wire[15:0] addr_selector3_2915;
wire[15:0] addr_remain3_2915;
address_decode_4 decoder_3_2915 = address_decode_4(addr_selector2_182[3],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2915,addr_remain3_2915);


wire[15:0] addr_selector3_2916;
wire[15:0] addr_remain3_2916;
address_decode_4 decoder_3_2916 = address_decode_4(addr_selector2_182[4],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2916,addr_remain3_2916);


wire[15:0] addr_selector3_2917;
wire[15:0] addr_remain3_2917;
address_decode_4 decoder_3_2917 = address_decode_4(addr_selector2_182[5],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2917,addr_remain3_2917);


wire[15:0] addr_selector3_2918;
wire[15:0] addr_remain3_2918;
address_decode_4 decoder_3_2918 = address_decode_4(addr_selector2_182[6],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2918,addr_remain3_2918);


wire[15:0] addr_selector3_2919;
wire[15:0] addr_remain3_2919;
address_decode_4 decoder_3_2919 = address_decode_4(addr_selector2_182[7],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2919,addr_remain3_2919);


wire[15:0] addr_selector3_2920;
wire[15:0] addr_remain3_2920;
address_decode_4 decoder_3_2920 = address_decode_4(addr_selector2_182[8],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2920,addr_remain3_2920);


wire[15:0] addr_selector3_2921;
wire[15:0] addr_remain3_2921;
address_decode_4 decoder_3_2921 = address_decode_4(addr_selector2_182[9],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2921,addr_remain3_2921);


wire[15:0] addr_selector3_2922;
wire[15:0] addr_remain3_2922;
address_decode_4 decoder_3_2922 = address_decode_4(addr_selector2_182[10],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2922,addr_remain3_2922);


wire[15:0] addr_selector3_2923;
wire[15:0] addr_remain3_2923;
address_decode_4 decoder_3_2923 = address_decode_4(addr_selector2_182[11],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2923,addr_remain3_2923);


wire[15:0] addr_selector3_2924;
wire[15:0] addr_remain3_2924;
address_decode_4 decoder_3_2924 = address_decode_4(addr_selector2_182[12],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2924,addr_remain3_2924);


wire[15:0] addr_selector3_2925;
wire[15:0] addr_remain3_2925;
address_decode_4 decoder_3_2925 = address_decode_4(addr_selector2_182[13],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2925,addr_remain3_2925);


wire[15:0] addr_selector3_2926;
wire[15:0] addr_remain3_2926;
address_decode_4 decoder_3_2926 = address_decode_4(addr_selector2_182[14],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2926,addr_remain3_2926);


wire[15:0] addr_selector3_2927;
wire[15:0] addr_remain3_2927;
address_decode_4 decoder_3_2927 = address_decode_4(addr_selector2_182[15],addr_remain2_182[15:0],addr_remain2_182,addr_selector3_2927,addr_remain3_2927);


wire[15:0] addr_selector3_2928;
wire[15:0] addr_remain3_2928;
address_decode_4 decoder_3_2928 = address_decode_4(addr_selector2_183[0],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2928,addr_remain3_2928);


wire[15:0] addr_selector3_2929;
wire[15:0] addr_remain3_2929;
address_decode_4 decoder_3_2929 = address_decode_4(addr_selector2_183[1],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2929,addr_remain3_2929);


wire[15:0] addr_selector3_2930;
wire[15:0] addr_remain3_2930;
address_decode_4 decoder_3_2930 = address_decode_4(addr_selector2_183[2],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2930,addr_remain3_2930);


wire[15:0] addr_selector3_2931;
wire[15:0] addr_remain3_2931;
address_decode_4 decoder_3_2931 = address_decode_4(addr_selector2_183[3],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2931,addr_remain3_2931);


wire[15:0] addr_selector3_2932;
wire[15:0] addr_remain3_2932;
address_decode_4 decoder_3_2932 = address_decode_4(addr_selector2_183[4],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2932,addr_remain3_2932);


wire[15:0] addr_selector3_2933;
wire[15:0] addr_remain3_2933;
address_decode_4 decoder_3_2933 = address_decode_4(addr_selector2_183[5],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2933,addr_remain3_2933);


wire[15:0] addr_selector3_2934;
wire[15:0] addr_remain3_2934;
address_decode_4 decoder_3_2934 = address_decode_4(addr_selector2_183[6],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2934,addr_remain3_2934);


wire[15:0] addr_selector3_2935;
wire[15:0] addr_remain3_2935;
address_decode_4 decoder_3_2935 = address_decode_4(addr_selector2_183[7],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2935,addr_remain3_2935);


wire[15:0] addr_selector3_2936;
wire[15:0] addr_remain3_2936;
address_decode_4 decoder_3_2936 = address_decode_4(addr_selector2_183[8],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2936,addr_remain3_2936);


wire[15:0] addr_selector3_2937;
wire[15:0] addr_remain3_2937;
address_decode_4 decoder_3_2937 = address_decode_4(addr_selector2_183[9],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2937,addr_remain3_2937);


wire[15:0] addr_selector3_2938;
wire[15:0] addr_remain3_2938;
address_decode_4 decoder_3_2938 = address_decode_4(addr_selector2_183[10],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2938,addr_remain3_2938);


wire[15:0] addr_selector3_2939;
wire[15:0] addr_remain3_2939;
address_decode_4 decoder_3_2939 = address_decode_4(addr_selector2_183[11],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2939,addr_remain3_2939);


wire[15:0] addr_selector3_2940;
wire[15:0] addr_remain3_2940;
address_decode_4 decoder_3_2940 = address_decode_4(addr_selector2_183[12],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2940,addr_remain3_2940);


wire[15:0] addr_selector3_2941;
wire[15:0] addr_remain3_2941;
address_decode_4 decoder_3_2941 = address_decode_4(addr_selector2_183[13],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2941,addr_remain3_2941);


wire[15:0] addr_selector3_2942;
wire[15:0] addr_remain3_2942;
address_decode_4 decoder_3_2942 = address_decode_4(addr_selector2_183[14],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2942,addr_remain3_2942);


wire[15:0] addr_selector3_2943;
wire[15:0] addr_remain3_2943;
address_decode_4 decoder_3_2943 = address_decode_4(addr_selector2_183[15],addr_remain2_183[15:0],addr_remain2_183,addr_selector3_2943,addr_remain3_2943);


wire[15:0] addr_selector3_2944;
wire[15:0] addr_remain3_2944;
address_decode_4 decoder_3_2944 = address_decode_4(addr_selector2_184[0],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2944,addr_remain3_2944);


wire[15:0] addr_selector3_2945;
wire[15:0] addr_remain3_2945;
address_decode_4 decoder_3_2945 = address_decode_4(addr_selector2_184[1],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2945,addr_remain3_2945);


wire[15:0] addr_selector3_2946;
wire[15:0] addr_remain3_2946;
address_decode_4 decoder_3_2946 = address_decode_4(addr_selector2_184[2],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2946,addr_remain3_2946);


wire[15:0] addr_selector3_2947;
wire[15:0] addr_remain3_2947;
address_decode_4 decoder_3_2947 = address_decode_4(addr_selector2_184[3],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2947,addr_remain3_2947);


wire[15:0] addr_selector3_2948;
wire[15:0] addr_remain3_2948;
address_decode_4 decoder_3_2948 = address_decode_4(addr_selector2_184[4],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2948,addr_remain3_2948);


wire[15:0] addr_selector3_2949;
wire[15:0] addr_remain3_2949;
address_decode_4 decoder_3_2949 = address_decode_4(addr_selector2_184[5],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2949,addr_remain3_2949);


wire[15:0] addr_selector3_2950;
wire[15:0] addr_remain3_2950;
address_decode_4 decoder_3_2950 = address_decode_4(addr_selector2_184[6],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2950,addr_remain3_2950);


wire[15:0] addr_selector3_2951;
wire[15:0] addr_remain3_2951;
address_decode_4 decoder_3_2951 = address_decode_4(addr_selector2_184[7],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2951,addr_remain3_2951);


wire[15:0] addr_selector3_2952;
wire[15:0] addr_remain3_2952;
address_decode_4 decoder_3_2952 = address_decode_4(addr_selector2_184[8],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2952,addr_remain3_2952);


wire[15:0] addr_selector3_2953;
wire[15:0] addr_remain3_2953;
address_decode_4 decoder_3_2953 = address_decode_4(addr_selector2_184[9],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2953,addr_remain3_2953);


wire[15:0] addr_selector3_2954;
wire[15:0] addr_remain3_2954;
address_decode_4 decoder_3_2954 = address_decode_4(addr_selector2_184[10],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2954,addr_remain3_2954);


wire[15:0] addr_selector3_2955;
wire[15:0] addr_remain3_2955;
address_decode_4 decoder_3_2955 = address_decode_4(addr_selector2_184[11],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2955,addr_remain3_2955);


wire[15:0] addr_selector3_2956;
wire[15:0] addr_remain3_2956;
address_decode_4 decoder_3_2956 = address_decode_4(addr_selector2_184[12],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2956,addr_remain3_2956);


wire[15:0] addr_selector3_2957;
wire[15:0] addr_remain3_2957;
address_decode_4 decoder_3_2957 = address_decode_4(addr_selector2_184[13],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2957,addr_remain3_2957);


wire[15:0] addr_selector3_2958;
wire[15:0] addr_remain3_2958;
address_decode_4 decoder_3_2958 = address_decode_4(addr_selector2_184[14],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2958,addr_remain3_2958);


wire[15:0] addr_selector3_2959;
wire[15:0] addr_remain3_2959;
address_decode_4 decoder_3_2959 = address_decode_4(addr_selector2_184[15],addr_remain2_184[15:0],addr_remain2_184,addr_selector3_2959,addr_remain3_2959);


wire[15:0] addr_selector3_2960;
wire[15:0] addr_remain3_2960;
address_decode_4 decoder_3_2960 = address_decode_4(addr_selector2_185[0],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2960,addr_remain3_2960);


wire[15:0] addr_selector3_2961;
wire[15:0] addr_remain3_2961;
address_decode_4 decoder_3_2961 = address_decode_4(addr_selector2_185[1],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2961,addr_remain3_2961);


wire[15:0] addr_selector3_2962;
wire[15:0] addr_remain3_2962;
address_decode_4 decoder_3_2962 = address_decode_4(addr_selector2_185[2],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2962,addr_remain3_2962);


wire[15:0] addr_selector3_2963;
wire[15:0] addr_remain3_2963;
address_decode_4 decoder_3_2963 = address_decode_4(addr_selector2_185[3],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2963,addr_remain3_2963);


wire[15:0] addr_selector3_2964;
wire[15:0] addr_remain3_2964;
address_decode_4 decoder_3_2964 = address_decode_4(addr_selector2_185[4],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2964,addr_remain3_2964);


wire[15:0] addr_selector3_2965;
wire[15:0] addr_remain3_2965;
address_decode_4 decoder_3_2965 = address_decode_4(addr_selector2_185[5],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2965,addr_remain3_2965);


wire[15:0] addr_selector3_2966;
wire[15:0] addr_remain3_2966;
address_decode_4 decoder_3_2966 = address_decode_4(addr_selector2_185[6],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2966,addr_remain3_2966);


wire[15:0] addr_selector3_2967;
wire[15:0] addr_remain3_2967;
address_decode_4 decoder_3_2967 = address_decode_4(addr_selector2_185[7],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2967,addr_remain3_2967);


wire[15:0] addr_selector3_2968;
wire[15:0] addr_remain3_2968;
address_decode_4 decoder_3_2968 = address_decode_4(addr_selector2_185[8],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2968,addr_remain3_2968);


wire[15:0] addr_selector3_2969;
wire[15:0] addr_remain3_2969;
address_decode_4 decoder_3_2969 = address_decode_4(addr_selector2_185[9],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2969,addr_remain3_2969);


wire[15:0] addr_selector3_2970;
wire[15:0] addr_remain3_2970;
address_decode_4 decoder_3_2970 = address_decode_4(addr_selector2_185[10],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2970,addr_remain3_2970);


wire[15:0] addr_selector3_2971;
wire[15:0] addr_remain3_2971;
address_decode_4 decoder_3_2971 = address_decode_4(addr_selector2_185[11],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2971,addr_remain3_2971);


wire[15:0] addr_selector3_2972;
wire[15:0] addr_remain3_2972;
address_decode_4 decoder_3_2972 = address_decode_4(addr_selector2_185[12],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2972,addr_remain3_2972);


wire[15:0] addr_selector3_2973;
wire[15:0] addr_remain3_2973;
address_decode_4 decoder_3_2973 = address_decode_4(addr_selector2_185[13],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2973,addr_remain3_2973);


wire[15:0] addr_selector3_2974;
wire[15:0] addr_remain3_2974;
address_decode_4 decoder_3_2974 = address_decode_4(addr_selector2_185[14],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2974,addr_remain3_2974);


wire[15:0] addr_selector3_2975;
wire[15:0] addr_remain3_2975;
address_decode_4 decoder_3_2975 = address_decode_4(addr_selector2_185[15],addr_remain2_185[15:0],addr_remain2_185,addr_selector3_2975,addr_remain3_2975);


wire[15:0] addr_selector3_2976;
wire[15:0] addr_remain3_2976;
address_decode_4 decoder_3_2976 = address_decode_4(addr_selector2_186[0],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2976,addr_remain3_2976);


wire[15:0] addr_selector3_2977;
wire[15:0] addr_remain3_2977;
address_decode_4 decoder_3_2977 = address_decode_4(addr_selector2_186[1],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2977,addr_remain3_2977);


wire[15:0] addr_selector3_2978;
wire[15:0] addr_remain3_2978;
address_decode_4 decoder_3_2978 = address_decode_4(addr_selector2_186[2],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2978,addr_remain3_2978);


wire[15:0] addr_selector3_2979;
wire[15:0] addr_remain3_2979;
address_decode_4 decoder_3_2979 = address_decode_4(addr_selector2_186[3],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2979,addr_remain3_2979);


wire[15:0] addr_selector3_2980;
wire[15:0] addr_remain3_2980;
address_decode_4 decoder_3_2980 = address_decode_4(addr_selector2_186[4],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2980,addr_remain3_2980);


wire[15:0] addr_selector3_2981;
wire[15:0] addr_remain3_2981;
address_decode_4 decoder_3_2981 = address_decode_4(addr_selector2_186[5],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2981,addr_remain3_2981);


wire[15:0] addr_selector3_2982;
wire[15:0] addr_remain3_2982;
address_decode_4 decoder_3_2982 = address_decode_4(addr_selector2_186[6],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2982,addr_remain3_2982);


wire[15:0] addr_selector3_2983;
wire[15:0] addr_remain3_2983;
address_decode_4 decoder_3_2983 = address_decode_4(addr_selector2_186[7],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2983,addr_remain3_2983);


wire[15:0] addr_selector3_2984;
wire[15:0] addr_remain3_2984;
address_decode_4 decoder_3_2984 = address_decode_4(addr_selector2_186[8],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2984,addr_remain3_2984);


wire[15:0] addr_selector3_2985;
wire[15:0] addr_remain3_2985;
address_decode_4 decoder_3_2985 = address_decode_4(addr_selector2_186[9],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2985,addr_remain3_2985);


wire[15:0] addr_selector3_2986;
wire[15:0] addr_remain3_2986;
address_decode_4 decoder_3_2986 = address_decode_4(addr_selector2_186[10],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2986,addr_remain3_2986);


wire[15:0] addr_selector3_2987;
wire[15:0] addr_remain3_2987;
address_decode_4 decoder_3_2987 = address_decode_4(addr_selector2_186[11],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2987,addr_remain3_2987);


wire[15:0] addr_selector3_2988;
wire[15:0] addr_remain3_2988;
address_decode_4 decoder_3_2988 = address_decode_4(addr_selector2_186[12],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2988,addr_remain3_2988);


wire[15:0] addr_selector3_2989;
wire[15:0] addr_remain3_2989;
address_decode_4 decoder_3_2989 = address_decode_4(addr_selector2_186[13],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2989,addr_remain3_2989);


wire[15:0] addr_selector3_2990;
wire[15:0] addr_remain3_2990;
address_decode_4 decoder_3_2990 = address_decode_4(addr_selector2_186[14],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2990,addr_remain3_2990);


wire[15:0] addr_selector3_2991;
wire[15:0] addr_remain3_2991;
address_decode_4 decoder_3_2991 = address_decode_4(addr_selector2_186[15],addr_remain2_186[15:0],addr_remain2_186,addr_selector3_2991,addr_remain3_2991);


wire[15:0] addr_selector3_2992;
wire[15:0] addr_remain3_2992;
address_decode_4 decoder_3_2992 = address_decode_4(addr_selector2_187[0],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2992,addr_remain3_2992);


wire[15:0] addr_selector3_2993;
wire[15:0] addr_remain3_2993;
address_decode_4 decoder_3_2993 = address_decode_4(addr_selector2_187[1],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2993,addr_remain3_2993);


wire[15:0] addr_selector3_2994;
wire[15:0] addr_remain3_2994;
address_decode_4 decoder_3_2994 = address_decode_4(addr_selector2_187[2],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2994,addr_remain3_2994);


wire[15:0] addr_selector3_2995;
wire[15:0] addr_remain3_2995;
address_decode_4 decoder_3_2995 = address_decode_4(addr_selector2_187[3],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2995,addr_remain3_2995);


wire[15:0] addr_selector3_2996;
wire[15:0] addr_remain3_2996;
address_decode_4 decoder_3_2996 = address_decode_4(addr_selector2_187[4],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2996,addr_remain3_2996);


wire[15:0] addr_selector3_2997;
wire[15:0] addr_remain3_2997;
address_decode_4 decoder_3_2997 = address_decode_4(addr_selector2_187[5],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2997,addr_remain3_2997);


wire[15:0] addr_selector3_2998;
wire[15:0] addr_remain3_2998;
address_decode_4 decoder_3_2998 = address_decode_4(addr_selector2_187[6],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2998,addr_remain3_2998);


wire[15:0] addr_selector3_2999;
wire[15:0] addr_remain3_2999;
address_decode_4 decoder_3_2999 = address_decode_4(addr_selector2_187[7],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_2999,addr_remain3_2999);


wire[15:0] addr_selector3_3000;
wire[15:0] addr_remain3_3000;
address_decode_4 decoder_3_3000 = address_decode_4(addr_selector2_187[8],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3000,addr_remain3_3000);


wire[15:0] addr_selector3_3001;
wire[15:0] addr_remain3_3001;
address_decode_4 decoder_3_3001 = address_decode_4(addr_selector2_187[9],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3001,addr_remain3_3001);


wire[15:0] addr_selector3_3002;
wire[15:0] addr_remain3_3002;
address_decode_4 decoder_3_3002 = address_decode_4(addr_selector2_187[10],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3002,addr_remain3_3002);


wire[15:0] addr_selector3_3003;
wire[15:0] addr_remain3_3003;
address_decode_4 decoder_3_3003 = address_decode_4(addr_selector2_187[11],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3003,addr_remain3_3003);


wire[15:0] addr_selector3_3004;
wire[15:0] addr_remain3_3004;
address_decode_4 decoder_3_3004 = address_decode_4(addr_selector2_187[12],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3004,addr_remain3_3004);


wire[15:0] addr_selector3_3005;
wire[15:0] addr_remain3_3005;
address_decode_4 decoder_3_3005 = address_decode_4(addr_selector2_187[13],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3005,addr_remain3_3005);


wire[15:0] addr_selector3_3006;
wire[15:0] addr_remain3_3006;
address_decode_4 decoder_3_3006 = address_decode_4(addr_selector2_187[14],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3006,addr_remain3_3006);


wire[15:0] addr_selector3_3007;
wire[15:0] addr_remain3_3007;
address_decode_4 decoder_3_3007 = address_decode_4(addr_selector2_187[15],addr_remain2_187[15:0],addr_remain2_187,addr_selector3_3007,addr_remain3_3007);


wire[15:0] addr_selector3_3008;
wire[15:0] addr_remain3_3008;
address_decode_4 decoder_3_3008 = address_decode_4(addr_selector2_188[0],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3008,addr_remain3_3008);


wire[15:0] addr_selector3_3009;
wire[15:0] addr_remain3_3009;
address_decode_4 decoder_3_3009 = address_decode_4(addr_selector2_188[1],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3009,addr_remain3_3009);


wire[15:0] addr_selector3_3010;
wire[15:0] addr_remain3_3010;
address_decode_4 decoder_3_3010 = address_decode_4(addr_selector2_188[2],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3010,addr_remain3_3010);


wire[15:0] addr_selector3_3011;
wire[15:0] addr_remain3_3011;
address_decode_4 decoder_3_3011 = address_decode_4(addr_selector2_188[3],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3011,addr_remain3_3011);


wire[15:0] addr_selector3_3012;
wire[15:0] addr_remain3_3012;
address_decode_4 decoder_3_3012 = address_decode_4(addr_selector2_188[4],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3012,addr_remain3_3012);


wire[15:0] addr_selector3_3013;
wire[15:0] addr_remain3_3013;
address_decode_4 decoder_3_3013 = address_decode_4(addr_selector2_188[5],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3013,addr_remain3_3013);


wire[15:0] addr_selector3_3014;
wire[15:0] addr_remain3_3014;
address_decode_4 decoder_3_3014 = address_decode_4(addr_selector2_188[6],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3014,addr_remain3_3014);


wire[15:0] addr_selector3_3015;
wire[15:0] addr_remain3_3015;
address_decode_4 decoder_3_3015 = address_decode_4(addr_selector2_188[7],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3015,addr_remain3_3015);


wire[15:0] addr_selector3_3016;
wire[15:0] addr_remain3_3016;
address_decode_4 decoder_3_3016 = address_decode_4(addr_selector2_188[8],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3016,addr_remain3_3016);


wire[15:0] addr_selector3_3017;
wire[15:0] addr_remain3_3017;
address_decode_4 decoder_3_3017 = address_decode_4(addr_selector2_188[9],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3017,addr_remain3_3017);


wire[15:0] addr_selector3_3018;
wire[15:0] addr_remain3_3018;
address_decode_4 decoder_3_3018 = address_decode_4(addr_selector2_188[10],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3018,addr_remain3_3018);


wire[15:0] addr_selector3_3019;
wire[15:0] addr_remain3_3019;
address_decode_4 decoder_3_3019 = address_decode_4(addr_selector2_188[11],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3019,addr_remain3_3019);


wire[15:0] addr_selector3_3020;
wire[15:0] addr_remain3_3020;
address_decode_4 decoder_3_3020 = address_decode_4(addr_selector2_188[12],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3020,addr_remain3_3020);


wire[15:0] addr_selector3_3021;
wire[15:0] addr_remain3_3021;
address_decode_4 decoder_3_3021 = address_decode_4(addr_selector2_188[13],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3021,addr_remain3_3021);


wire[15:0] addr_selector3_3022;
wire[15:0] addr_remain3_3022;
address_decode_4 decoder_3_3022 = address_decode_4(addr_selector2_188[14],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3022,addr_remain3_3022);


wire[15:0] addr_selector3_3023;
wire[15:0] addr_remain3_3023;
address_decode_4 decoder_3_3023 = address_decode_4(addr_selector2_188[15],addr_remain2_188[15:0],addr_remain2_188,addr_selector3_3023,addr_remain3_3023);


wire[15:0] addr_selector3_3024;
wire[15:0] addr_remain3_3024;
address_decode_4 decoder_3_3024 = address_decode_4(addr_selector2_189[0],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3024,addr_remain3_3024);


wire[15:0] addr_selector3_3025;
wire[15:0] addr_remain3_3025;
address_decode_4 decoder_3_3025 = address_decode_4(addr_selector2_189[1],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3025,addr_remain3_3025);


wire[15:0] addr_selector3_3026;
wire[15:0] addr_remain3_3026;
address_decode_4 decoder_3_3026 = address_decode_4(addr_selector2_189[2],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3026,addr_remain3_3026);


wire[15:0] addr_selector3_3027;
wire[15:0] addr_remain3_3027;
address_decode_4 decoder_3_3027 = address_decode_4(addr_selector2_189[3],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3027,addr_remain3_3027);


wire[15:0] addr_selector3_3028;
wire[15:0] addr_remain3_3028;
address_decode_4 decoder_3_3028 = address_decode_4(addr_selector2_189[4],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3028,addr_remain3_3028);


wire[15:0] addr_selector3_3029;
wire[15:0] addr_remain3_3029;
address_decode_4 decoder_3_3029 = address_decode_4(addr_selector2_189[5],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3029,addr_remain3_3029);


wire[15:0] addr_selector3_3030;
wire[15:0] addr_remain3_3030;
address_decode_4 decoder_3_3030 = address_decode_4(addr_selector2_189[6],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3030,addr_remain3_3030);


wire[15:0] addr_selector3_3031;
wire[15:0] addr_remain3_3031;
address_decode_4 decoder_3_3031 = address_decode_4(addr_selector2_189[7],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3031,addr_remain3_3031);


wire[15:0] addr_selector3_3032;
wire[15:0] addr_remain3_3032;
address_decode_4 decoder_3_3032 = address_decode_4(addr_selector2_189[8],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3032,addr_remain3_3032);


wire[15:0] addr_selector3_3033;
wire[15:0] addr_remain3_3033;
address_decode_4 decoder_3_3033 = address_decode_4(addr_selector2_189[9],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3033,addr_remain3_3033);


wire[15:0] addr_selector3_3034;
wire[15:0] addr_remain3_3034;
address_decode_4 decoder_3_3034 = address_decode_4(addr_selector2_189[10],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3034,addr_remain3_3034);


wire[15:0] addr_selector3_3035;
wire[15:0] addr_remain3_3035;
address_decode_4 decoder_3_3035 = address_decode_4(addr_selector2_189[11],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3035,addr_remain3_3035);


wire[15:0] addr_selector3_3036;
wire[15:0] addr_remain3_3036;
address_decode_4 decoder_3_3036 = address_decode_4(addr_selector2_189[12],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3036,addr_remain3_3036);


wire[15:0] addr_selector3_3037;
wire[15:0] addr_remain3_3037;
address_decode_4 decoder_3_3037 = address_decode_4(addr_selector2_189[13],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3037,addr_remain3_3037);


wire[15:0] addr_selector3_3038;
wire[15:0] addr_remain3_3038;
address_decode_4 decoder_3_3038 = address_decode_4(addr_selector2_189[14],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3038,addr_remain3_3038);


wire[15:0] addr_selector3_3039;
wire[15:0] addr_remain3_3039;
address_decode_4 decoder_3_3039 = address_decode_4(addr_selector2_189[15],addr_remain2_189[15:0],addr_remain2_189,addr_selector3_3039,addr_remain3_3039);


wire[15:0] addr_selector3_3040;
wire[15:0] addr_remain3_3040;
address_decode_4 decoder_3_3040 = address_decode_4(addr_selector2_190[0],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3040,addr_remain3_3040);


wire[15:0] addr_selector3_3041;
wire[15:0] addr_remain3_3041;
address_decode_4 decoder_3_3041 = address_decode_4(addr_selector2_190[1],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3041,addr_remain3_3041);


wire[15:0] addr_selector3_3042;
wire[15:0] addr_remain3_3042;
address_decode_4 decoder_3_3042 = address_decode_4(addr_selector2_190[2],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3042,addr_remain3_3042);


wire[15:0] addr_selector3_3043;
wire[15:0] addr_remain3_3043;
address_decode_4 decoder_3_3043 = address_decode_4(addr_selector2_190[3],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3043,addr_remain3_3043);


wire[15:0] addr_selector3_3044;
wire[15:0] addr_remain3_3044;
address_decode_4 decoder_3_3044 = address_decode_4(addr_selector2_190[4],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3044,addr_remain3_3044);


wire[15:0] addr_selector3_3045;
wire[15:0] addr_remain3_3045;
address_decode_4 decoder_3_3045 = address_decode_4(addr_selector2_190[5],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3045,addr_remain3_3045);


wire[15:0] addr_selector3_3046;
wire[15:0] addr_remain3_3046;
address_decode_4 decoder_3_3046 = address_decode_4(addr_selector2_190[6],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3046,addr_remain3_3046);


wire[15:0] addr_selector3_3047;
wire[15:0] addr_remain3_3047;
address_decode_4 decoder_3_3047 = address_decode_4(addr_selector2_190[7],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3047,addr_remain3_3047);


wire[15:0] addr_selector3_3048;
wire[15:0] addr_remain3_3048;
address_decode_4 decoder_3_3048 = address_decode_4(addr_selector2_190[8],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3048,addr_remain3_3048);


wire[15:0] addr_selector3_3049;
wire[15:0] addr_remain3_3049;
address_decode_4 decoder_3_3049 = address_decode_4(addr_selector2_190[9],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3049,addr_remain3_3049);


wire[15:0] addr_selector3_3050;
wire[15:0] addr_remain3_3050;
address_decode_4 decoder_3_3050 = address_decode_4(addr_selector2_190[10],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3050,addr_remain3_3050);


wire[15:0] addr_selector3_3051;
wire[15:0] addr_remain3_3051;
address_decode_4 decoder_3_3051 = address_decode_4(addr_selector2_190[11],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3051,addr_remain3_3051);


wire[15:0] addr_selector3_3052;
wire[15:0] addr_remain3_3052;
address_decode_4 decoder_3_3052 = address_decode_4(addr_selector2_190[12],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3052,addr_remain3_3052);


wire[15:0] addr_selector3_3053;
wire[15:0] addr_remain3_3053;
address_decode_4 decoder_3_3053 = address_decode_4(addr_selector2_190[13],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3053,addr_remain3_3053);


wire[15:0] addr_selector3_3054;
wire[15:0] addr_remain3_3054;
address_decode_4 decoder_3_3054 = address_decode_4(addr_selector2_190[14],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3054,addr_remain3_3054);


wire[15:0] addr_selector3_3055;
wire[15:0] addr_remain3_3055;
address_decode_4 decoder_3_3055 = address_decode_4(addr_selector2_190[15],addr_remain2_190[15:0],addr_remain2_190,addr_selector3_3055,addr_remain3_3055);


wire[15:0] addr_selector3_3056;
wire[15:0] addr_remain3_3056;
address_decode_4 decoder_3_3056 = address_decode_4(addr_selector2_191[0],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3056,addr_remain3_3056);


wire[15:0] addr_selector3_3057;
wire[15:0] addr_remain3_3057;
address_decode_4 decoder_3_3057 = address_decode_4(addr_selector2_191[1],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3057,addr_remain3_3057);


wire[15:0] addr_selector3_3058;
wire[15:0] addr_remain3_3058;
address_decode_4 decoder_3_3058 = address_decode_4(addr_selector2_191[2],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3058,addr_remain3_3058);


wire[15:0] addr_selector3_3059;
wire[15:0] addr_remain3_3059;
address_decode_4 decoder_3_3059 = address_decode_4(addr_selector2_191[3],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3059,addr_remain3_3059);


wire[15:0] addr_selector3_3060;
wire[15:0] addr_remain3_3060;
address_decode_4 decoder_3_3060 = address_decode_4(addr_selector2_191[4],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3060,addr_remain3_3060);


wire[15:0] addr_selector3_3061;
wire[15:0] addr_remain3_3061;
address_decode_4 decoder_3_3061 = address_decode_4(addr_selector2_191[5],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3061,addr_remain3_3061);


wire[15:0] addr_selector3_3062;
wire[15:0] addr_remain3_3062;
address_decode_4 decoder_3_3062 = address_decode_4(addr_selector2_191[6],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3062,addr_remain3_3062);


wire[15:0] addr_selector3_3063;
wire[15:0] addr_remain3_3063;
address_decode_4 decoder_3_3063 = address_decode_4(addr_selector2_191[7],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3063,addr_remain3_3063);


wire[15:0] addr_selector3_3064;
wire[15:0] addr_remain3_3064;
address_decode_4 decoder_3_3064 = address_decode_4(addr_selector2_191[8],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3064,addr_remain3_3064);


wire[15:0] addr_selector3_3065;
wire[15:0] addr_remain3_3065;
address_decode_4 decoder_3_3065 = address_decode_4(addr_selector2_191[9],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3065,addr_remain3_3065);


wire[15:0] addr_selector3_3066;
wire[15:0] addr_remain3_3066;
address_decode_4 decoder_3_3066 = address_decode_4(addr_selector2_191[10],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3066,addr_remain3_3066);


wire[15:0] addr_selector3_3067;
wire[15:0] addr_remain3_3067;
address_decode_4 decoder_3_3067 = address_decode_4(addr_selector2_191[11],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3067,addr_remain3_3067);


wire[15:0] addr_selector3_3068;
wire[15:0] addr_remain3_3068;
address_decode_4 decoder_3_3068 = address_decode_4(addr_selector2_191[12],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3068,addr_remain3_3068);


wire[15:0] addr_selector3_3069;
wire[15:0] addr_remain3_3069;
address_decode_4 decoder_3_3069 = address_decode_4(addr_selector2_191[13],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3069,addr_remain3_3069);


wire[15:0] addr_selector3_3070;
wire[15:0] addr_remain3_3070;
address_decode_4 decoder_3_3070 = address_decode_4(addr_selector2_191[14],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3070,addr_remain3_3070);


wire[15:0] addr_selector3_3071;
wire[15:0] addr_remain3_3071;
address_decode_4 decoder_3_3071 = address_decode_4(addr_selector2_191[15],addr_remain2_191[15:0],addr_remain2_191,addr_selector3_3071,addr_remain3_3071);


wire[15:0] addr_selector3_3072;
wire[15:0] addr_remain3_3072;
address_decode_4 decoder_3_3072 = address_decode_4(addr_selector2_192[0],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3072,addr_remain3_3072);


wire[15:0] addr_selector3_3073;
wire[15:0] addr_remain3_3073;
address_decode_4 decoder_3_3073 = address_decode_4(addr_selector2_192[1],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3073,addr_remain3_3073);


wire[15:0] addr_selector3_3074;
wire[15:0] addr_remain3_3074;
address_decode_4 decoder_3_3074 = address_decode_4(addr_selector2_192[2],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3074,addr_remain3_3074);


wire[15:0] addr_selector3_3075;
wire[15:0] addr_remain3_3075;
address_decode_4 decoder_3_3075 = address_decode_4(addr_selector2_192[3],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3075,addr_remain3_3075);


wire[15:0] addr_selector3_3076;
wire[15:0] addr_remain3_3076;
address_decode_4 decoder_3_3076 = address_decode_4(addr_selector2_192[4],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3076,addr_remain3_3076);


wire[15:0] addr_selector3_3077;
wire[15:0] addr_remain3_3077;
address_decode_4 decoder_3_3077 = address_decode_4(addr_selector2_192[5],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3077,addr_remain3_3077);


wire[15:0] addr_selector3_3078;
wire[15:0] addr_remain3_3078;
address_decode_4 decoder_3_3078 = address_decode_4(addr_selector2_192[6],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3078,addr_remain3_3078);


wire[15:0] addr_selector3_3079;
wire[15:0] addr_remain3_3079;
address_decode_4 decoder_3_3079 = address_decode_4(addr_selector2_192[7],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3079,addr_remain3_3079);


wire[15:0] addr_selector3_3080;
wire[15:0] addr_remain3_3080;
address_decode_4 decoder_3_3080 = address_decode_4(addr_selector2_192[8],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3080,addr_remain3_3080);


wire[15:0] addr_selector3_3081;
wire[15:0] addr_remain3_3081;
address_decode_4 decoder_3_3081 = address_decode_4(addr_selector2_192[9],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3081,addr_remain3_3081);


wire[15:0] addr_selector3_3082;
wire[15:0] addr_remain3_3082;
address_decode_4 decoder_3_3082 = address_decode_4(addr_selector2_192[10],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3082,addr_remain3_3082);


wire[15:0] addr_selector3_3083;
wire[15:0] addr_remain3_3083;
address_decode_4 decoder_3_3083 = address_decode_4(addr_selector2_192[11],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3083,addr_remain3_3083);


wire[15:0] addr_selector3_3084;
wire[15:0] addr_remain3_3084;
address_decode_4 decoder_3_3084 = address_decode_4(addr_selector2_192[12],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3084,addr_remain3_3084);


wire[15:0] addr_selector3_3085;
wire[15:0] addr_remain3_3085;
address_decode_4 decoder_3_3085 = address_decode_4(addr_selector2_192[13],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3085,addr_remain3_3085);


wire[15:0] addr_selector3_3086;
wire[15:0] addr_remain3_3086;
address_decode_4 decoder_3_3086 = address_decode_4(addr_selector2_192[14],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3086,addr_remain3_3086);


wire[15:0] addr_selector3_3087;
wire[15:0] addr_remain3_3087;
address_decode_4 decoder_3_3087 = address_decode_4(addr_selector2_192[15],addr_remain2_192[15:0],addr_remain2_192,addr_selector3_3087,addr_remain3_3087);


wire[15:0] addr_selector3_3088;
wire[15:0] addr_remain3_3088;
address_decode_4 decoder_3_3088 = address_decode_4(addr_selector2_193[0],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3088,addr_remain3_3088);


wire[15:0] addr_selector3_3089;
wire[15:0] addr_remain3_3089;
address_decode_4 decoder_3_3089 = address_decode_4(addr_selector2_193[1],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3089,addr_remain3_3089);


wire[15:0] addr_selector3_3090;
wire[15:0] addr_remain3_3090;
address_decode_4 decoder_3_3090 = address_decode_4(addr_selector2_193[2],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3090,addr_remain3_3090);


wire[15:0] addr_selector3_3091;
wire[15:0] addr_remain3_3091;
address_decode_4 decoder_3_3091 = address_decode_4(addr_selector2_193[3],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3091,addr_remain3_3091);


wire[15:0] addr_selector3_3092;
wire[15:0] addr_remain3_3092;
address_decode_4 decoder_3_3092 = address_decode_4(addr_selector2_193[4],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3092,addr_remain3_3092);


wire[15:0] addr_selector3_3093;
wire[15:0] addr_remain3_3093;
address_decode_4 decoder_3_3093 = address_decode_4(addr_selector2_193[5],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3093,addr_remain3_3093);


wire[15:0] addr_selector3_3094;
wire[15:0] addr_remain3_3094;
address_decode_4 decoder_3_3094 = address_decode_4(addr_selector2_193[6],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3094,addr_remain3_3094);


wire[15:0] addr_selector3_3095;
wire[15:0] addr_remain3_3095;
address_decode_4 decoder_3_3095 = address_decode_4(addr_selector2_193[7],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3095,addr_remain3_3095);


wire[15:0] addr_selector3_3096;
wire[15:0] addr_remain3_3096;
address_decode_4 decoder_3_3096 = address_decode_4(addr_selector2_193[8],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3096,addr_remain3_3096);


wire[15:0] addr_selector3_3097;
wire[15:0] addr_remain3_3097;
address_decode_4 decoder_3_3097 = address_decode_4(addr_selector2_193[9],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3097,addr_remain3_3097);


wire[15:0] addr_selector3_3098;
wire[15:0] addr_remain3_3098;
address_decode_4 decoder_3_3098 = address_decode_4(addr_selector2_193[10],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3098,addr_remain3_3098);


wire[15:0] addr_selector3_3099;
wire[15:0] addr_remain3_3099;
address_decode_4 decoder_3_3099 = address_decode_4(addr_selector2_193[11],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3099,addr_remain3_3099);


wire[15:0] addr_selector3_3100;
wire[15:0] addr_remain3_3100;
address_decode_4 decoder_3_3100 = address_decode_4(addr_selector2_193[12],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3100,addr_remain3_3100);


wire[15:0] addr_selector3_3101;
wire[15:0] addr_remain3_3101;
address_decode_4 decoder_3_3101 = address_decode_4(addr_selector2_193[13],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3101,addr_remain3_3101);


wire[15:0] addr_selector3_3102;
wire[15:0] addr_remain3_3102;
address_decode_4 decoder_3_3102 = address_decode_4(addr_selector2_193[14],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3102,addr_remain3_3102);


wire[15:0] addr_selector3_3103;
wire[15:0] addr_remain3_3103;
address_decode_4 decoder_3_3103 = address_decode_4(addr_selector2_193[15],addr_remain2_193[15:0],addr_remain2_193,addr_selector3_3103,addr_remain3_3103);


wire[15:0] addr_selector3_3104;
wire[15:0] addr_remain3_3104;
address_decode_4 decoder_3_3104 = address_decode_4(addr_selector2_194[0],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3104,addr_remain3_3104);


wire[15:0] addr_selector3_3105;
wire[15:0] addr_remain3_3105;
address_decode_4 decoder_3_3105 = address_decode_4(addr_selector2_194[1],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3105,addr_remain3_3105);


wire[15:0] addr_selector3_3106;
wire[15:0] addr_remain3_3106;
address_decode_4 decoder_3_3106 = address_decode_4(addr_selector2_194[2],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3106,addr_remain3_3106);


wire[15:0] addr_selector3_3107;
wire[15:0] addr_remain3_3107;
address_decode_4 decoder_3_3107 = address_decode_4(addr_selector2_194[3],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3107,addr_remain3_3107);


wire[15:0] addr_selector3_3108;
wire[15:0] addr_remain3_3108;
address_decode_4 decoder_3_3108 = address_decode_4(addr_selector2_194[4],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3108,addr_remain3_3108);


wire[15:0] addr_selector3_3109;
wire[15:0] addr_remain3_3109;
address_decode_4 decoder_3_3109 = address_decode_4(addr_selector2_194[5],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3109,addr_remain3_3109);


wire[15:0] addr_selector3_3110;
wire[15:0] addr_remain3_3110;
address_decode_4 decoder_3_3110 = address_decode_4(addr_selector2_194[6],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3110,addr_remain3_3110);


wire[15:0] addr_selector3_3111;
wire[15:0] addr_remain3_3111;
address_decode_4 decoder_3_3111 = address_decode_4(addr_selector2_194[7],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3111,addr_remain3_3111);


wire[15:0] addr_selector3_3112;
wire[15:0] addr_remain3_3112;
address_decode_4 decoder_3_3112 = address_decode_4(addr_selector2_194[8],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3112,addr_remain3_3112);


wire[15:0] addr_selector3_3113;
wire[15:0] addr_remain3_3113;
address_decode_4 decoder_3_3113 = address_decode_4(addr_selector2_194[9],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3113,addr_remain3_3113);


wire[15:0] addr_selector3_3114;
wire[15:0] addr_remain3_3114;
address_decode_4 decoder_3_3114 = address_decode_4(addr_selector2_194[10],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3114,addr_remain3_3114);


wire[15:0] addr_selector3_3115;
wire[15:0] addr_remain3_3115;
address_decode_4 decoder_3_3115 = address_decode_4(addr_selector2_194[11],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3115,addr_remain3_3115);


wire[15:0] addr_selector3_3116;
wire[15:0] addr_remain3_3116;
address_decode_4 decoder_3_3116 = address_decode_4(addr_selector2_194[12],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3116,addr_remain3_3116);


wire[15:0] addr_selector3_3117;
wire[15:0] addr_remain3_3117;
address_decode_4 decoder_3_3117 = address_decode_4(addr_selector2_194[13],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3117,addr_remain3_3117);


wire[15:0] addr_selector3_3118;
wire[15:0] addr_remain3_3118;
address_decode_4 decoder_3_3118 = address_decode_4(addr_selector2_194[14],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3118,addr_remain3_3118);


wire[15:0] addr_selector3_3119;
wire[15:0] addr_remain3_3119;
address_decode_4 decoder_3_3119 = address_decode_4(addr_selector2_194[15],addr_remain2_194[15:0],addr_remain2_194,addr_selector3_3119,addr_remain3_3119);


wire[15:0] addr_selector3_3120;
wire[15:0] addr_remain3_3120;
address_decode_4 decoder_3_3120 = address_decode_4(addr_selector2_195[0],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3120,addr_remain3_3120);


wire[15:0] addr_selector3_3121;
wire[15:0] addr_remain3_3121;
address_decode_4 decoder_3_3121 = address_decode_4(addr_selector2_195[1],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3121,addr_remain3_3121);


wire[15:0] addr_selector3_3122;
wire[15:0] addr_remain3_3122;
address_decode_4 decoder_3_3122 = address_decode_4(addr_selector2_195[2],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3122,addr_remain3_3122);


wire[15:0] addr_selector3_3123;
wire[15:0] addr_remain3_3123;
address_decode_4 decoder_3_3123 = address_decode_4(addr_selector2_195[3],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3123,addr_remain3_3123);


wire[15:0] addr_selector3_3124;
wire[15:0] addr_remain3_3124;
address_decode_4 decoder_3_3124 = address_decode_4(addr_selector2_195[4],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3124,addr_remain3_3124);


wire[15:0] addr_selector3_3125;
wire[15:0] addr_remain3_3125;
address_decode_4 decoder_3_3125 = address_decode_4(addr_selector2_195[5],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3125,addr_remain3_3125);


wire[15:0] addr_selector3_3126;
wire[15:0] addr_remain3_3126;
address_decode_4 decoder_3_3126 = address_decode_4(addr_selector2_195[6],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3126,addr_remain3_3126);


wire[15:0] addr_selector3_3127;
wire[15:0] addr_remain3_3127;
address_decode_4 decoder_3_3127 = address_decode_4(addr_selector2_195[7],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3127,addr_remain3_3127);


wire[15:0] addr_selector3_3128;
wire[15:0] addr_remain3_3128;
address_decode_4 decoder_3_3128 = address_decode_4(addr_selector2_195[8],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3128,addr_remain3_3128);


wire[15:0] addr_selector3_3129;
wire[15:0] addr_remain3_3129;
address_decode_4 decoder_3_3129 = address_decode_4(addr_selector2_195[9],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3129,addr_remain3_3129);


wire[15:0] addr_selector3_3130;
wire[15:0] addr_remain3_3130;
address_decode_4 decoder_3_3130 = address_decode_4(addr_selector2_195[10],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3130,addr_remain3_3130);


wire[15:0] addr_selector3_3131;
wire[15:0] addr_remain3_3131;
address_decode_4 decoder_3_3131 = address_decode_4(addr_selector2_195[11],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3131,addr_remain3_3131);


wire[15:0] addr_selector3_3132;
wire[15:0] addr_remain3_3132;
address_decode_4 decoder_3_3132 = address_decode_4(addr_selector2_195[12],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3132,addr_remain3_3132);


wire[15:0] addr_selector3_3133;
wire[15:0] addr_remain3_3133;
address_decode_4 decoder_3_3133 = address_decode_4(addr_selector2_195[13],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3133,addr_remain3_3133);


wire[15:0] addr_selector3_3134;
wire[15:0] addr_remain3_3134;
address_decode_4 decoder_3_3134 = address_decode_4(addr_selector2_195[14],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3134,addr_remain3_3134);


wire[15:0] addr_selector3_3135;
wire[15:0] addr_remain3_3135;
address_decode_4 decoder_3_3135 = address_decode_4(addr_selector2_195[15],addr_remain2_195[15:0],addr_remain2_195,addr_selector3_3135,addr_remain3_3135);


wire[15:0] addr_selector3_3136;
wire[15:0] addr_remain3_3136;
address_decode_4 decoder_3_3136 = address_decode_4(addr_selector2_196[0],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3136,addr_remain3_3136);


wire[15:0] addr_selector3_3137;
wire[15:0] addr_remain3_3137;
address_decode_4 decoder_3_3137 = address_decode_4(addr_selector2_196[1],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3137,addr_remain3_3137);


wire[15:0] addr_selector3_3138;
wire[15:0] addr_remain3_3138;
address_decode_4 decoder_3_3138 = address_decode_4(addr_selector2_196[2],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3138,addr_remain3_3138);


wire[15:0] addr_selector3_3139;
wire[15:0] addr_remain3_3139;
address_decode_4 decoder_3_3139 = address_decode_4(addr_selector2_196[3],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3139,addr_remain3_3139);


wire[15:0] addr_selector3_3140;
wire[15:0] addr_remain3_3140;
address_decode_4 decoder_3_3140 = address_decode_4(addr_selector2_196[4],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3140,addr_remain3_3140);


wire[15:0] addr_selector3_3141;
wire[15:0] addr_remain3_3141;
address_decode_4 decoder_3_3141 = address_decode_4(addr_selector2_196[5],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3141,addr_remain3_3141);


wire[15:0] addr_selector3_3142;
wire[15:0] addr_remain3_3142;
address_decode_4 decoder_3_3142 = address_decode_4(addr_selector2_196[6],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3142,addr_remain3_3142);


wire[15:0] addr_selector3_3143;
wire[15:0] addr_remain3_3143;
address_decode_4 decoder_3_3143 = address_decode_4(addr_selector2_196[7],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3143,addr_remain3_3143);


wire[15:0] addr_selector3_3144;
wire[15:0] addr_remain3_3144;
address_decode_4 decoder_3_3144 = address_decode_4(addr_selector2_196[8],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3144,addr_remain3_3144);


wire[15:0] addr_selector3_3145;
wire[15:0] addr_remain3_3145;
address_decode_4 decoder_3_3145 = address_decode_4(addr_selector2_196[9],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3145,addr_remain3_3145);


wire[15:0] addr_selector3_3146;
wire[15:0] addr_remain3_3146;
address_decode_4 decoder_3_3146 = address_decode_4(addr_selector2_196[10],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3146,addr_remain3_3146);


wire[15:0] addr_selector3_3147;
wire[15:0] addr_remain3_3147;
address_decode_4 decoder_3_3147 = address_decode_4(addr_selector2_196[11],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3147,addr_remain3_3147);


wire[15:0] addr_selector3_3148;
wire[15:0] addr_remain3_3148;
address_decode_4 decoder_3_3148 = address_decode_4(addr_selector2_196[12],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3148,addr_remain3_3148);


wire[15:0] addr_selector3_3149;
wire[15:0] addr_remain3_3149;
address_decode_4 decoder_3_3149 = address_decode_4(addr_selector2_196[13],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3149,addr_remain3_3149);


wire[15:0] addr_selector3_3150;
wire[15:0] addr_remain3_3150;
address_decode_4 decoder_3_3150 = address_decode_4(addr_selector2_196[14],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3150,addr_remain3_3150);


wire[15:0] addr_selector3_3151;
wire[15:0] addr_remain3_3151;
address_decode_4 decoder_3_3151 = address_decode_4(addr_selector2_196[15],addr_remain2_196[15:0],addr_remain2_196,addr_selector3_3151,addr_remain3_3151);


wire[15:0] addr_selector3_3152;
wire[15:0] addr_remain3_3152;
address_decode_4 decoder_3_3152 = address_decode_4(addr_selector2_197[0],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3152,addr_remain3_3152);


wire[15:0] addr_selector3_3153;
wire[15:0] addr_remain3_3153;
address_decode_4 decoder_3_3153 = address_decode_4(addr_selector2_197[1],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3153,addr_remain3_3153);


wire[15:0] addr_selector3_3154;
wire[15:0] addr_remain3_3154;
address_decode_4 decoder_3_3154 = address_decode_4(addr_selector2_197[2],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3154,addr_remain3_3154);


wire[15:0] addr_selector3_3155;
wire[15:0] addr_remain3_3155;
address_decode_4 decoder_3_3155 = address_decode_4(addr_selector2_197[3],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3155,addr_remain3_3155);


wire[15:0] addr_selector3_3156;
wire[15:0] addr_remain3_3156;
address_decode_4 decoder_3_3156 = address_decode_4(addr_selector2_197[4],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3156,addr_remain3_3156);


wire[15:0] addr_selector3_3157;
wire[15:0] addr_remain3_3157;
address_decode_4 decoder_3_3157 = address_decode_4(addr_selector2_197[5],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3157,addr_remain3_3157);


wire[15:0] addr_selector3_3158;
wire[15:0] addr_remain3_3158;
address_decode_4 decoder_3_3158 = address_decode_4(addr_selector2_197[6],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3158,addr_remain3_3158);


wire[15:0] addr_selector3_3159;
wire[15:0] addr_remain3_3159;
address_decode_4 decoder_3_3159 = address_decode_4(addr_selector2_197[7],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3159,addr_remain3_3159);


wire[15:0] addr_selector3_3160;
wire[15:0] addr_remain3_3160;
address_decode_4 decoder_3_3160 = address_decode_4(addr_selector2_197[8],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3160,addr_remain3_3160);


wire[15:0] addr_selector3_3161;
wire[15:0] addr_remain3_3161;
address_decode_4 decoder_3_3161 = address_decode_4(addr_selector2_197[9],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3161,addr_remain3_3161);


wire[15:0] addr_selector3_3162;
wire[15:0] addr_remain3_3162;
address_decode_4 decoder_3_3162 = address_decode_4(addr_selector2_197[10],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3162,addr_remain3_3162);


wire[15:0] addr_selector3_3163;
wire[15:0] addr_remain3_3163;
address_decode_4 decoder_3_3163 = address_decode_4(addr_selector2_197[11],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3163,addr_remain3_3163);


wire[15:0] addr_selector3_3164;
wire[15:0] addr_remain3_3164;
address_decode_4 decoder_3_3164 = address_decode_4(addr_selector2_197[12],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3164,addr_remain3_3164);


wire[15:0] addr_selector3_3165;
wire[15:0] addr_remain3_3165;
address_decode_4 decoder_3_3165 = address_decode_4(addr_selector2_197[13],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3165,addr_remain3_3165);


wire[15:0] addr_selector3_3166;
wire[15:0] addr_remain3_3166;
address_decode_4 decoder_3_3166 = address_decode_4(addr_selector2_197[14],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3166,addr_remain3_3166);


wire[15:0] addr_selector3_3167;
wire[15:0] addr_remain3_3167;
address_decode_4 decoder_3_3167 = address_decode_4(addr_selector2_197[15],addr_remain2_197[15:0],addr_remain2_197,addr_selector3_3167,addr_remain3_3167);


wire[15:0] addr_selector3_3168;
wire[15:0] addr_remain3_3168;
address_decode_4 decoder_3_3168 = address_decode_4(addr_selector2_198[0],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3168,addr_remain3_3168);


wire[15:0] addr_selector3_3169;
wire[15:0] addr_remain3_3169;
address_decode_4 decoder_3_3169 = address_decode_4(addr_selector2_198[1],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3169,addr_remain3_3169);


wire[15:0] addr_selector3_3170;
wire[15:0] addr_remain3_3170;
address_decode_4 decoder_3_3170 = address_decode_4(addr_selector2_198[2],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3170,addr_remain3_3170);


wire[15:0] addr_selector3_3171;
wire[15:0] addr_remain3_3171;
address_decode_4 decoder_3_3171 = address_decode_4(addr_selector2_198[3],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3171,addr_remain3_3171);


wire[15:0] addr_selector3_3172;
wire[15:0] addr_remain3_3172;
address_decode_4 decoder_3_3172 = address_decode_4(addr_selector2_198[4],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3172,addr_remain3_3172);


wire[15:0] addr_selector3_3173;
wire[15:0] addr_remain3_3173;
address_decode_4 decoder_3_3173 = address_decode_4(addr_selector2_198[5],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3173,addr_remain3_3173);


wire[15:0] addr_selector3_3174;
wire[15:0] addr_remain3_3174;
address_decode_4 decoder_3_3174 = address_decode_4(addr_selector2_198[6],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3174,addr_remain3_3174);


wire[15:0] addr_selector3_3175;
wire[15:0] addr_remain3_3175;
address_decode_4 decoder_3_3175 = address_decode_4(addr_selector2_198[7],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3175,addr_remain3_3175);


wire[15:0] addr_selector3_3176;
wire[15:0] addr_remain3_3176;
address_decode_4 decoder_3_3176 = address_decode_4(addr_selector2_198[8],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3176,addr_remain3_3176);


wire[15:0] addr_selector3_3177;
wire[15:0] addr_remain3_3177;
address_decode_4 decoder_3_3177 = address_decode_4(addr_selector2_198[9],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3177,addr_remain3_3177);


wire[15:0] addr_selector3_3178;
wire[15:0] addr_remain3_3178;
address_decode_4 decoder_3_3178 = address_decode_4(addr_selector2_198[10],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3178,addr_remain3_3178);


wire[15:0] addr_selector3_3179;
wire[15:0] addr_remain3_3179;
address_decode_4 decoder_3_3179 = address_decode_4(addr_selector2_198[11],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3179,addr_remain3_3179);


wire[15:0] addr_selector3_3180;
wire[15:0] addr_remain3_3180;
address_decode_4 decoder_3_3180 = address_decode_4(addr_selector2_198[12],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3180,addr_remain3_3180);


wire[15:0] addr_selector3_3181;
wire[15:0] addr_remain3_3181;
address_decode_4 decoder_3_3181 = address_decode_4(addr_selector2_198[13],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3181,addr_remain3_3181);


wire[15:0] addr_selector3_3182;
wire[15:0] addr_remain3_3182;
address_decode_4 decoder_3_3182 = address_decode_4(addr_selector2_198[14],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3182,addr_remain3_3182);


wire[15:0] addr_selector3_3183;
wire[15:0] addr_remain3_3183;
address_decode_4 decoder_3_3183 = address_decode_4(addr_selector2_198[15],addr_remain2_198[15:0],addr_remain2_198,addr_selector3_3183,addr_remain3_3183);


wire[15:0] addr_selector3_3184;
wire[15:0] addr_remain3_3184;
address_decode_4 decoder_3_3184 = address_decode_4(addr_selector2_199[0],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3184,addr_remain3_3184);


wire[15:0] addr_selector3_3185;
wire[15:0] addr_remain3_3185;
address_decode_4 decoder_3_3185 = address_decode_4(addr_selector2_199[1],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3185,addr_remain3_3185);


wire[15:0] addr_selector3_3186;
wire[15:0] addr_remain3_3186;
address_decode_4 decoder_3_3186 = address_decode_4(addr_selector2_199[2],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3186,addr_remain3_3186);


wire[15:0] addr_selector3_3187;
wire[15:0] addr_remain3_3187;
address_decode_4 decoder_3_3187 = address_decode_4(addr_selector2_199[3],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3187,addr_remain3_3187);


wire[15:0] addr_selector3_3188;
wire[15:0] addr_remain3_3188;
address_decode_4 decoder_3_3188 = address_decode_4(addr_selector2_199[4],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3188,addr_remain3_3188);


wire[15:0] addr_selector3_3189;
wire[15:0] addr_remain3_3189;
address_decode_4 decoder_3_3189 = address_decode_4(addr_selector2_199[5],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3189,addr_remain3_3189);


wire[15:0] addr_selector3_3190;
wire[15:0] addr_remain3_3190;
address_decode_4 decoder_3_3190 = address_decode_4(addr_selector2_199[6],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3190,addr_remain3_3190);


wire[15:0] addr_selector3_3191;
wire[15:0] addr_remain3_3191;
address_decode_4 decoder_3_3191 = address_decode_4(addr_selector2_199[7],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3191,addr_remain3_3191);


wire[15:0] addr_selector3_3192;
wire[15:0] addr_remain3_3192;
address_decode_4 decoder_3_3192 = address_decode_4(addr_selector2_199[8],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3192,addr_remain3_3192);


wire[15:0] addr_selector3_3193;
wire[15:0] addr_remain3_3193;
address_decode_4 decoder_3_3193 = address_decode_4(addr_selector2_199[9],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3193,addr_remain3_3193);


wire[15:0] addr_selector3_3194;
wire[15:0] addr_remain3_3194;
address_decode_4 decoder_3_3194 = address_decode_4(addr_selector2_199[10],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3194,addr_remain3_3194);


wire[15:0] addr_selector3_3195;
wire[15:0] addr_remain3_3195;
address_decode_4 decoder_3_3195 = address_decode_4(addr_selector2_199[11],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3195,addr_remain3_3195);


wire[15:0] addr_selector3_3196;
wire[15:0] addr_remain3_3196;
address_decode_4 decoder_3_3196 = address_decode_4(addr_selector2_199[12],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3196,addr_remain3_3196);


wire[15:0] addr_selector3_3197;
wire[15:0] addr_remain3_3197;
address_decode_4 decoder_3_3197 = address_decode_4(addr_selector2_199[13],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3197,addr_remain3_3197);


wire[15:0] addr_selector3_3198;
wire[15:0] addr_remain3_3198;
address_decode_4 decoder_3_3198 = address_decode_4(addr_selector2_199[14],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3198,addr_remain3_3198);


wire[15:0] addr_selector3_3199;
wire[15:0] addr_remain3_3199;
address_decode_4 decoder_3_3199 = address_decode_4(addr_selector2_199[15],addr_remain2_199[15:0],addr_remain2_199,addr_selector3_3199,addr_remain3_3199);


wire[15:0] addr_selector3_3200;
wire[15:0] addr_remain3_3200;
address_decode_4 decoder_3_3200 = address_decode_4(addr_selector2_200[0],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3200,addr_remain3_3200);


wire[15:0] addr_selector3_3201;
wire[15:0] addr_remain3_3201;
address_decode_4 decoder_3_3201 = address_decode_4(addr_selector2_200[1],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3201,addr_remain3_3201);


wire[15:0] addr_selector3_3202;
wire[15:0] addr_remain3_3202;
address_decode_4 decoder_3_3202 = address_decode_4(addr_selector2_200[2],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3202,addr_remain3_3202);


wire[15:0] addr_selector3_3203;
wire[15:0] addr_remain3_3203;
address_decode_4 decoder_3_3203 = address_decode_4(addr_selector2_200[3],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3203,addr_remain3_3203);


wire[15:0] addr_selector3_3204;
wire[15:0] addr_remain3_3204;
address_decode_4 decoder_3_3204 = address_decode_4(addr_selector2_200[4],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3204,addr_remain3_3204);


wire[15:0] addr_selector3_3205;
wire[15:0] addr_remain3_3205;
address_decode_4 decoder_3_3205 = address_decode_4(addr_selector2_200[5],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3205,addr_remain3_3205);


wire[15:0] addr_selector3_3206;
wire[15:0] addr_remain3_3206;
address_decode_4 decoder_3_3206 = address_decode_4(addr_selector2_200[6],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3206,addr_remain3_3206);


wire[15:0] addr_selector3_3207;
wire[15:0] addr_remain3_3207;
address_decode_4 decoder_3_3207 = address_decode_4(addr_selector2_200[7],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3207,addr_remain3_3207);


wire[15:0] addr_selector3_3208;
wire[15:0] addr_remain3_3208;
address_decode_4 decoder_3_3208 = address_decode_4(addr_selector2_200[8],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3208,addr_remain3_3208);


wire[15:0] addr_selector3_3209;
wire[15:0] addr_remain3_3209;
address_decode_4 decoder_3_3209 = address_decode_4(addr_selector2_200[9],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3209,addr_remain3_3209);


wire[15:0] addr_selector3_3210;
wire[15:0] addr_remain3_3210;
address_decode_4 decoder_3_3210 = address_decode_4(addr_selector2_200[10],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3210,addr_remain3_3210);


wire[15:0] addr_selector3_3211;
wire[15:0] addr_remain3_3211;
address_decode_4 decoder_3_3211 = address_decode_4(addr_selector2_200[11],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3211,addr_remain3_3211);


wire[15:0] addr_selector3_3212;
wire[15:0] addr_remain3_3212;
address_decode_4 decoder_3_3212 = address_decode_4(addr_selector2_200[12],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3212,addr_remain3_3212);


wire[15:0] addr_selector3_3213;
wire[15:0] addr_remain3_3213;
address_decode_4 decoder_3_3213 = address_decode_4(addr_selector2_200[13],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3213,addr_remain3_3213);


wire[15:0] addr_selector3_3214;
wire[15:0] addr_remain3_3214;
address_decode_4 decoder_3_3214 = address_decode_4(addr_selector2_200[14],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3214,addr_remain3_3214);


wire[15:0] addr_selector3_3215;
wire[15:0] addr_remain3_3215;
address_decode_4 decoder_3_3215 = address_decode_4(addr_selector2_200[15],addr_remain2_200[15:0],addr_remain2_200,addr_selector3_3215,addr_remain3_3215);


wire[15:0] addr_selector3_3216;
wire[15:0] addr_remain3_3216;
address_decode_4 decoder_3_3216 = address_decode_4(addr_selector2_201[0],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3216,addr_remain3_3216);


wire[15:0] addr_selector3_3217;
wire[15:0] addr_remain3_3217;
address_decode_4 decoder_3_3217 = address_decode_4(addr_selector2_201[1],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3217,addr_remain3_3217);


wire[15:0] addr_selector3_3218;
wire[15:0] addr_remain3_3218;
address_decode_4 decoder_3_3218 = address_decode_4(addr_selector2_201[2],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3218,addr_remain3_3218);


wire[15:0] addr_selector3_3219;
wire[15:0] addr_remain3_3219;
address_decode_4 decoder_3_3219 = address_decode_4(addr_selector2_201[3],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3219,addr_remain3_3219);


wire[15:0] addr_selector3_3220;
wire[15:0] addr_remain3_3220;
address_decode_4 decoder_3_3220 = address_decode_4(addr_selector2_201[4],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3220,addr_remain3_3220);


wire[15:0] addr_selector3_3221;
wire[15:0] addr_remain3_3221;
address_decode_4 decoder_3_3221 = address_decode_4(addr_selector2_201[5],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3221,addr_remain3_3221);


wire[15:0] addr_selector3_3222;
wire[15:0] addr_remain3_3222;
address_decode_4 decoder_3_3222 = address_decode_4(addr_selector2_201[6],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3222,addr_remain3_3222);


wire[15:0] addr_selector3_3223;
wire[15:0] addr_remain3_3223;
address_decode_4 decoder_3_3223 = address_decode_4(addr_selector2_201[7],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3223,addr_remain3_3223);


wire[15:0] addr_selector3_3224;
wire[15:0] addr_remain3_3224;
address_decode_4 decoder_3_3224 = address_decode_4(addr_selector2_201[8],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3224,addr_remain3_3224);


wire[15:0] addr_selector3_3225;
wire[15:0] addr_remain3_3225;
address_decode_4 decoder_3_3225 = address_decode_4(addr_selector2_201[9],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3225,addr_remain3_3225);


wire[15:0] addr_selector3_3226;
wire[15:0] addr_remain3_3226;
address_decode_4 decoder_3_3226 = address_decode_4(addr_selector2_201[10],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3226,addr_remain3_3226);


wire[15:0] addr_selector3_3227;
wire[15:0] addr_remain3_3227;
address_decode_4 decoder_3_3227 = address_decode_4(addr_selector2_201[11],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3227,addr_remain3_3227);


wire[15:0] addr_selector3_3228;
wire[15:0] addr_remain3_3228;
address_decode_4 decoder_3_3228 = address_decode_4(addr_selector2_201[12],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3228,addr_remain3_3228);


wire[15:0] addr_selector3_3229;
wire[15:0] addr_remain3_3229;
address_decode_4 decoder_3_3229 = address_decode_4(addr_selector2_201[13],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3229,addr_remain3_3229);


wire[15:0] addr_selector3_3230;
wire[15:0] addr_remain3_3230;
address_decode_4 decoder_3_3230 = address_decode_4(addr_selector2_201[14],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3230,addr_remain3_3230);


wire[15:0] addr_selector3_3231;
wire[15:0] addr_remain3_3231;
address_decode_4 decoder_3_3231 = address_decode_4(addr_selector2_201[15],addr_remain2_201[15:0],addr_remain2_201,addr_selector3_3231,addr_remain3_3231);


wire[15:0] addr_selector3_3232;
wire[15:0] addr_remain3_3232;
address_decode_4 decoder_3_3232 = address_decode_4(addr_selector2_202[0],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3232,addr_remain3_3232);


wire[15:0] addr_selector3_3233;
wire[15:0] addr_remain3_3233;
address_decode_4 decoder_3_3233 = address_decode_4(addr_selector2_202[1],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3233,addr_remain3_3233);


wire[15:0] addr_selector3_3234;
wire[15:0] addr_remain3_3234;
address_decode_4 decoder_3_3234 = address_decode_4(addr_selector2_202[2],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3234,addr_remain3_3234);


wire[15:0] addr_selector3_3235;
wire[15:0] addr_remain3_3235;
address_decode_4 decoder_3_3235 = address_decode_4(addr_selector2_202[3],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3235,addr_remain3_3235);


wire[15:0] addr_selector3_3236;
wire[15:0] addr_remain3_3236;
address_decode_4 decoder_3_3236 = address_decode_4(addr_selector2_202[4],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3236,addr_remain3_3236);


wire[15:0] addr_selector3_3237;
wire[15:0] addr_remain3_3237;
address_decode_4 decoder_3_3237 = address_decode_4(addr_selector2_202[5],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3237,addr_remain3_3237);


wire[15:0] addr_selector3_3238;
wire[15:0] addr_remain3_3238;
address_decode_4 decoder_3_3238 = address_decode_4(addr_selector2_202[6],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3238,addr_remain3_3238);


wire[15:0] addr_selector3_3239;
wire[15:0] addr_remain3_3239;
address_decode_4 decoder_3_3239 = address_decode_4(addr_selector2_202[7],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3239,addr_remain3_3239);


wire[15:0] addr_selector3_3240;
wire[15:0] addr_remain3_3240;
address_decode_4 decoder_3_3240 = address_decode_4(addr_selector2_202[8],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3240,addr_remain3_3240);


wire[15:0] addr_selector3_3241;
wire[15:0] addr_remain3_3241;
address_decode_4 decoder_3_3241 = address_decode_4(addr_selector2_202[9],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3241,addr_remain3_3241);


wire[15:0] addr_selector3_3242;
wire[15:0] addr_remain3_3242;
address_decode_4 decoder_3_3242 = address_decode_4(addr_selector2_202[10],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3242,addr_remain3_3242);


wire[15:0] addr_selector3_3243;
wire[15:0] addr_remain3_3243;
address_decode_4 decoder_3_3243 = address_decode_4(addr_selector2_202[11],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3243,addr_remain3_3243);


wire[15:0] addr_selector3_3244;
wire[15:0] addr_remain3_3244;
address_decode_4 decoder_3_3244 = address_decode_4(addr_selector2_202[12],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3244,addr_remain3_3244);


wire[15:0] addr_selector3_3245;
wire[15:0] addr_remain3_3245;
address_decode_4 decoder_3_3245 = address_decode_4(addr_selector2_202[13],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3245,addr_remain3_3245);


wire[15:0] addr_selector3_3246;
wire[15:0] addr_remain3_3246;
address_decode_4 decoder_3_3246 = address_decode_4(addr_selector2_202[14],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3246,addr_remain3_3246);


wire[15:0] addr_selector3_3247;
wire[15:0] addr_remain3_3247;
address_decode_4 decoder_3_3247 = address_decode_4(addr_selector2_202[15],addr_remain2_202[15:0],addr_remain2_202,addr_selector3_3247,addr_remain3_3247);


wire[15:0] addr_selector3_3248;
wire[15:0] addr_remain3_3248;
address_decode_4 decoder_3_3248 = address_decode_4(addr_selector2_203[0],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3248,addr_remain3_3248);


wire[15:0] addr_selector3_3249;
wire[15:0] addr_remain3_3249;
address_decode_4 decoder_3_3249 = address_decode_4(addr_selector2_203[1],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3249,addr_remain3_3249);


wire[15:0] addr_selector3_3250;
wire[15:0] addr_remain3_3250;
address_decode_4 decoder_3_3250 = address_decode_4(addr_selector2_203[2],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3250,addr_remain3_3250);


wire[15:0] addr_selector3_3251;
wire[15:0] addr_remain3_3251;
address_decode_4 decoder_3_3251 = address_decode_4(addr_selector2_203[3],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3251,addr_remain3_3251);


wire[15:0] addr_selector3_3252;
wire[15:0] addr_remain3_3252;
address_decode_4 decoder_3_3252 = address_decode_4(addr_selector2_203[4],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3252,addr_remain3_3252);


wire[15:0] addr_selector3_3253;
wire[15:0] addr_remain3_3253;
address_decode_4 decoder_3_3253 = address_decode_4(addr_selector2_203[5],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3253,addr_remain3_3253);


wire[15:0] addr_selector3_3254;
wire[15:0] addr_remain3_3254;
address_decode_4 decoder_3_3254 = address_decode_4(addr_selector2_203[6],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3254,addr_remain3_3254);


wire[15:0] addr_selector3_3255;
wire[15:0] addr_remain3_3255;
address_decode_4 decoder_3_3255 = address_decode_4(addr_selector2_203[7],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3255,addr_remain3_3255);


wire[15:0] addr_selector3_3256;
wire[15:0] addr_remain3_3256;
address_decode_4 decoder_3_3256 = address_decode_4(addr_selector2_203[8],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3256,addr_remain3_3256);


wire[15:0] addr_selector3_3257;
wire[15:0] addr_remain3_3257;
address_decode_4 decoder_3_3257 = address_decode_4(addr_selector2_203[9],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3257,addr_remain3_3257);


wire[15:0] addr_selector3_3258;
wire[15:0] addr_remain3_3258;
address_decode_4 decoder_3_3258 = address_decode_4(addr_selector2_203[10],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3258,addr_remain3_3258);


wire[15:0] addr_selector3_3259;
wire[15:0] addr_remain3_3259;
address_decode_4 decoder_3_3259 = address_decode_4(addr_selector2_203[11],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3259,addr_remain3_3259);


wire[15:0] addr_selector3_3260;
wire[15:0] addr_remain3_3260;
address_decode_4 decoder_3_3260 = address_decode_4(addr_selector2_203[12],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3260,addr_remain3_3260);


wire[15:0] addr_selector3_3261;
wire[15:0] addr_remain3_3261;
address_decode_4 decoder_3_3261 = address_decode_4(addr_selector2_203[13],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3261,addr_remain3_3261);


wire[15:0] addr_selector3_3262;
wire[15:0] addr_remain3_3262;
address_decode_4 decoder_3_3262 = address_decode_4(addr_selector2_203[14],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3262,addr_remain3_3262);


wire[15:0] addr_selector3_3263;
wire[15:0] addr_remain3_3263;
address_decode_4 decoder_3_3263 = address_decode_4(addr_selector2_203[15],addr_remain2_203[15:0],addr_remain2_203,addr_selector3_3263,addr_remain3_3263);


wire[15:0] addr_selector3_3264;
wire[15:0] addr_remain3_3264;
address_decode_4 decoder_3_3264 = address_decode_4(addr_selector2_204[0],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3264,addr_remain3_3264);


wire[15:0] addr_selector3_3265;
wire[15:0] addr_remain3_3265;
address_decode_4 decoder_3_3265 = address_decode_4(addr_selector2_204[1],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3265,addr_remain3_3265);


wire[15:0] addr_selector3_3266;
wire[15:0] addr_remain3_3266;
address_decode_4 decoder_3_3266 = address_decode_4(addr_selector2_204[2],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3266,addr_remain3_3266);


wire[15:0] addr_selector3_3267;
wire[15:0] addr_remain3_3267;
address_decode_4 decoder_3_3267 = address_decode_4(addr_selector2_204[3],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3267,addr_remain3_3267);


wire[15:0] addr_selector3_3268;
wire[15:0] addr_remain3_3268;
address_decode_4 decoder_3_3268 = address_decode_4(addr_selector2_204[4],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3268,addr_remain3_3268);


wire[15:0] addr_selector3_3269;
wire[15:0] addr_remain3_3269;
address_decode_4 decoder_3_3269 = address_decode_4(addr_selector2_204[5],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3269,addr_remain3_3269);


wire[15:0] addr_selector3_3270;
wire[15:0] addr_remain3_3270;
address_decode_4 decoder_3_3270 = address_decode_4(addr_selector2_204[6],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3270,addr_remain3_3270);


wire[15:0] addr_selector3_3271;
wire[15:0] addr_remain3_3271;
address_decode_4 decoder_3_3271 = address_decode_4(addr_selector2_204[7],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3271,addr_remain3_3271);


wire[15:0] addr_selector3_3272;
wire[15:0] addr_remain3_3272;
address_decode_4 decoder_3_3272 = address_decode_4(addr_selector2_204[8],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3272,addr_remain3_3272);


wire[15:0] addr_selector3_3273;
wire[15:0] addr_remain3_3273;
address_decode_4 decoder_3_3273 = address_decode_4(addr_selector2_204[9],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3273,addr_remain3_3273);


wire[15:0] addr_selector3_3274;
wire[15:0] addr_remain3_3274;
address_decode_4 decoder_3_3274 = address_decode_4(addr_selector2_204[10],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3274,addr_remain3_3274);


wire[15:0] addr_selector3_3275;
wire[15:0] addr_remain3_3275;
address_decode_4 decoder_3_3275 = address_decode_4(addr_selector2_204[11],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3275,addr_remain3_3275);


wire[15:0] addr_selector3_3276;
wire[15:0] addr_remain3_3276;
address_decode_4 decoder_3_3276 = address_decode_4(addr_selector2_204[12],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3276,addr_remain3_3276);


wire[15:0] addr_selector3_3277;
wire[15:0] addr_remain3_3277;
address_decode_4 decoder_3_3277 = address_decode_4(addr_selector2_204[13],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3277,addr_remain3_3277);


wire[15:0] addr_selector3_3278;
wire[15:0] addr_remain3_3278;
address_decode_4 decoder_3_3278 = address_decode_4(addr_selector2_204[14],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3278,addr_remain3_3278);


wire[15:0] addr_selector3_3279;
wire[15:0] addr_remain3_3279;
address_decode_4 decoder_3_3279 = address_decode_4(addr_selector2_204[15],addr_remain2_204[15:0],addr_remain2_204,addr_selector3_3279,addr_remain3_3279);


wire[15:0] addr_selector3_3280;
wire[15:0] addr_remain3_3280;
address_decode_4 decoder_3_3280 = address_decode_4(addr_selector2_205[0],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3280,addr_remain3_3280);


wire[15:0] addr_selector3_3281;
wire[15:0] addr_remain3_3281;
address_decode_4 decoder_3_3281 = address_decode_4(addr_selector2_205[1],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3281,addr_remain3_3281);


wire[15:0] addr_selector3_3282;
wire[15:0] addr_remain3_3282;
address_decode_4 decoder_3_3282 = address_decode_4(addr_selector2_205[2],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3282,addr_remain3_3282);


wire[15:0] addr_selector3_3283;
wire[15:0] addr_remain3_3283;
address_decode_4 decoder_3_3283 = address_decode_4(addr_selector2_205[3],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3283,addr_remain3_3283);


wire[15:0] addr_selector3_3284;
wire[15:0] addr_remain3_3284;
address_decode_4 decoder_3_3284 = address_decode_4(addr_selector2_205[4],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3284,addr_remain3_3284);


wire[15:0] addr_selector3_3285;
wire[15:0] addr_remain3_3285;
address_decode_4 decoder_3_3285 = address_decode_4(addr_selector2_205[5],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3285,addr_remain3_3285);


wire[15:0] addr_selector3_3286;
wire[15:0] addr_remain3_3286;
address_decode_4 decoder_3_3286 = address_decode_4(addr_selector2_205[6],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3286,addr_remain3_3286);


wire[15:0] addr_selector3_3287;
wire[15:0] addr_remain3_3287;
address_decode_4 decoder_3_3287 = address_decode_4(addr_selector2_205[7],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3287,addr_remain3_3287);


wire[15:0] addr_selector3_3288;
wire[15:0] addr_remain3_3288;
address_decode_4 decoder_3_3288 = address_decode_4(addr_selector2_205[8],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3288,addr_remain3_3288);


wire[15:0] addr_selector3_3289;
wire[15:0] addr_remain3_3289;
address_decode_4 decoder_3_3289 = address_decode_4(addr_selector2_205[9],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3289,addr_remain3_3289);


wire[15:0] addr_selector3_3290;
wire[15:0] addr_remain3_3290;
address_decode_4 decoder_3_3290 = address_decode_4(addr_selector2_205[10],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3290,addr_remain3_3290);


wire[15:0] addr_selector3_3291;
wire[15:0] addr_remain3_3291;
address_decode_4 decoder_3_3291 = address_decode_4(addr_selector2_205[11],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3291,addr_remain3_3291);


wire[15:0] addr_selector3_3292;
wire[15:0] addr_remain3_3292;
address_decode_4 decoder_3_3292 = address_decode_4(addr_selector2_205[12],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3292,addr_remain3_3292);


wire[15:0] addr_selector3_3293;
wire[15:0] addr_remain3_3293;
address_decode_4 decoder_3_3293 = address_decode_4(addr_selector2_205[13],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3293,addr_remain3_3293);


wire[15:0] addr_selector3_3294;
wire[15:0] addr_remain3_3294;
address_decode_4 decoder_3_3294 = address_decode_4(addr_selector2_205[14],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3294,addr_remain3_3294);


wire[15:0] addr_selector3_3295;
wire[15:0] addr_remain3_3295;
address_decode_4 decoder_3_3295 = address_decode_4(addr_selector2_205[15],addr_remain2_205[15:0],addr_remain2_205,addr_selector3_3295,addr_remain3_3295);


wire[15:0] addr_selector3_3296;
wire[15:0] addr_remain3_3296;
address_decode_4 decoder_3_3296 = address_decode_4(addr_selector2_206[0],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3296,addr_remain3_3296);


wire[15:0] addr_selector3_3297;
wire[15:0] addr_remain3_3297;
address_decode_4 decoder_3_3297 = address_decode_4(addr_selector2_206[1],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3297,addr_remain3_3297);


wire[15:0] addr_selector3_3298;
wire[15:0] addr_remain3_3298;
address_decode_4 decoder_3_3298 = address_decode_4(addr_selector2_206[2],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3298,addr_remain3_3298);


wire[15:0] addr_selector3_3299;
wire[15:0] addr_remain3_3299;
address_decode_4 decoder_3_3299 = address_decode_4(addr_selector2_206[3],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3299,addr_remain3_3299);


wire[15:0] addr_selector3_3300;
wire[15:0] addr_remain3_3300;
address_decode_4 decoder_3_3300 = address_decode_4(addr_selector2_206[4],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3300,addr_remain3_3300);


wire[15:0] addr_selector3_3301;
wire[15:0] addr_remain3_3301;
address_decode_4 decoder_3_3301 = address_decode_4(addr_selector2_206[5],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3301,addr_remain3_3301);


wire[15:0] addr_selector3_3302;
wire[15:0] addr_remain3_3302;
address_decode_4 decoder_3_3302 = address_decode_4(addr_selector2_206[6],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3302,addr_remain3_3302);


wire[15:0] addr_selector3_3303;
wire[15:0] addr_remain3_3303;
address_decode_4 decoder_3_3303 = address_decode_4(addr_selector2_206[7],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3303,addr_remain3_3303);


wire[15:0] addr_selector3_3304;
wire[15:0] addr_remain3_3304;
address_decode_4 decoder_3_3304 = address_decode_4(addr_selector2_206[8],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3304,addr_remain3_3304);


wire[15:0] addr_selector3_3305;
wire[15:0] addr_remain3_3305;
address_decode_4 decoder_3_3305 = address_decode_4(addr_selector2_206[9],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3305,addr_remain3_3305);


wire[15:0] addr_selector3_3306;
wire[15:0] addr_remain3_3306;
address_decode_4 decoder_3_3306 = address_decode_4(addr_selector2_206[10],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3306,addr_remain3_3306);


wire[15:0] addr_selector3_3307;
wire[15:0] addr_remain3_3307;
address_decode_4 decoder_3_3307 = address_decode_4(addr_selector2_206[11],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3307,addr_remain3_3307);


wire[15:0] addr_selector3_3308;
wire[15:0] addr_remain3_3308;
address_decode_4 decoder_3_3308 = address_decode_4(addr_selector2_206[12],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3308,addr_remain3_3308);


wire[15:0] addr_selector3_3309;
wire[15:0] addr_remain3_3309;
address_decode_4 decoder_3_3309 = address_decode_4(addr_selector2_206[13],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3309,addr_remain3_3309);


wire[15:0] addr_selector3_3310;
wire[15:0] addr_remain3_3310;
address_decode_4 decoder_3_3310 = address_decode_4(addr_selector2_206[14],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3310,addr_remain3_3310);


wire[15:0] addr_selector3_3311;
wire[15:0] addr_remain3_3311;
address_decode_4 decoder_3_3311 = address_decode_4(addr_selector2_206[15],addr_remain2_206[15:0],addr_remain2_206,addr_selector3_3311,addr_remain3_3311);


wire[15:0] addr_selector3_3312;
wire[15:0] addr_remain3_3312;
address_decode_4 decoder_3_3312 = address_decode_4(addr_selector2_207[0],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3312,addr_remain3_3312);


wire[15:0] addr_selector3_3313;
wire[15:0] addr_remain3_3313;
address_decode_4 decoder_3_3313 = address_decode_4(addr_selector2_207[1],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3313,addr_remain3_3313);


wire[15:0] addr_selector3_3314;
wire[15:0] addr_remain3_3314;
address_decode_4 decoder_3_3314 = address_decode_4(addr_selector2_207[2],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3314,addr_remain3_3314);


wire[15:0] addr_selector3_3315;
wire[15:0] addr_remain3_3315;
address_decode_4 decoder_3_3315 = address_decode_4(addr_selector2_207[3],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3315,addr_remain3_3315);


wire[15:0] addr_selector3_3316;
wire[15:0] addr_remain3_3316;
address_decode_4 decoder_3_3316 = address_decode_4(addr_selector2_207[4],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3316,addr_remain3_3316);


wire[15:0] addr_selector3_3317;
wire[15:0] addr_remain3_3317;
address_decode_4 decoder_3_3317 = address_decode_4(addr_selector2_207[5],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3317,addr_remain3_3317);


wire[15:0] addr_selector3_3318;
wire[15:0] addr_remain3_3318;
address_decode_4 decoder_3_3318 = address_decode_4(addr_selector2_207[6],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3318,addr_remain3_3318);


wire[15:0] addr_selector3_3319;
wire[15:0] addr_remain3_3319;
address_decode_4 decoder_3_3319 = address_decode_4(addr_selector2_207[7],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3319,addr_remain3_3319);


wire[15:0] addr_selector3_3320;
wire[15:0] addr_remain3_3320;
address_decode_4 decoder_3_3320 = address_decode_4(addr_selector2_207[8],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3320,addr_remain3_3320);


wire[15:0] addr_selector3_3321;
wire[15:0] addr_remain3_3321;
address_decode_4 decoder_3_3321 = address_decode_4(addr_selector2_207[9],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3321,addr_remain3_3321);


wire[15:0] addr_selector3_3322;
wire[15:0] addr_remain3_3322;
address_decode_4 decoder_3_3322 = address_decode_4(addr_selector2_207[10],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3322,addr_remain3_3322);


wire[15:0] addr_selector3_3323;
wire[15:0] addr_remain3_3323;
address_decode_4 decoder_3_3323 = address_decode_4(addr_selector2_207[11],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3323,addr_remain3_3323);


wire[15:0] addr_selector3_3324;
wire[15:0] addr_remain3_3324;
address_decode_4 decoder_3_3324 = address_decode_4(addr_selector2_207[12],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3324,addr_remain3_3324);


wire[15:0] addr_selector3_3325;
wire[15:0] addr_remain3_3325;
address_decode_4 decoder_3_3325 = address_decode_4(addr_selector2_207[13],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3325,addr_remain3_3325);


wire[15:0] addr_selector3_3326;
wire[15:0] addr_remain3_3326;
address_decode_4 decoder_3_3326 = address_decode_4(addr_selector2_207[14],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3326,addr_remain3_3326);


wire[15:0] addr_selector3_3327;
wire[15:0] addr_remain3_3327;
address_decode_4 decoder_3_3327 = address_decode_4(addr_selector2_207[15],addr_remain2_207[15:0],addr_remain2_207,addr_selector3_3327,addr_remain3_3327);


wire[15:0] addr_selector3_3328;
wire[15:0] addr_remain3_3328;
address_decode_4 decoder_3_3328 = address_decode_4(addr_selector2_208[0],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3328,addr_remain3_3328);


wire[15:0] addr_selector3_3329;
wire[15:0] addr_remain3_3329;
address_decode_4 decoder_3_3329 = address_decode_4(addr_selector2_208[1],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3329,addr_remain3_3329);


wire[15:0] addr_selector3_3330;
wire[15:0] addr_remain3_3330;
address_decode_4 decoder_3_3330 = address_decode_4(addr_selector2_208[2],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3330,addr_remain3_3330);


wire[15:0] addr_selector3_3331;
wire[15:0] addr_remain3_3331;
address_decode_4 decoder_3_3331 = address_decode_4(addr_selector2_208[3],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3331,addr_remain3_3331);


wire[15:0] addr_selector3_3332;
wire[15:0] addr_remain3_3332;
address_decode_4 decoder_3_3332 = address_decode_4(addr_selector2_208[4],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3332,addr_remain3_3332);


wire[15:0] addr_selector3_3333;
wire[15:0] addr_remain3_3333;
address_decode_4 decoder_3_3333 = address_decode_4(addr_selector2_208[5],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3333,addr_remain3_3333);


wire[15:0] addr_selector3_3334;
wire[15:0] addr_remain3_3334;
address_decode_4 decoder_3_3334 = address_decode_4(addr_selector2_208[6],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3334,addr_remain3_3334);


wire[15:0] addr_selector3_3335;
wire[15:0] addr_remain3_3335;
address_decode_4 decoder_3_3335 = address_decode_4(addr_selector2_208[7],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3335,addr_remain3_3335);


wire[15:0] addr_selector3_3336;
wire[15:0] addr_remain3_3336;
address_decode_4 decoder_3_3336 = address_decode_4(addr_selector2_208[8],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3336,addr_remain3_3336);


wire[15:0] addr_selector3_3337;
wire[15:0] addr_remain3_3337;
address_decode_4 decoder_3_3337 = address_decode_4(addr_selector2_208[9],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3337,addr_remain3_3337);


wire[15:0] addr_selector3_3338;
wire[15:0] addr_remain3_3338;
address_decode_4 decoder_3_3338 = address_decode_4(addr_selector2_208[10],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3338,addr_remain3_3338);


wire[15:0] addr_selector3_3339;
wire[15:0] addr_remain3_3339;
address_decode_4 decoder_3_3339 = address_decode_4(addr_selector2_208[11],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3339,addr_remain3_3339);


wire[15:0] addr_selector3_3340;
wire[15:0] addr_remain3_3340;
address_decode_4 decoder_3_3340 = address_decode_4(addr_selector2_208[12],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3340,addr_remain3_3340);


wire[15:0] addr_selector3_3341;
wire[15:0] addr_remain3_3341;
address_decode_4 decoder_3_3341 = address_decode_4(addr_selector2_208[13],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3341,addr_remain3_3341);


wire[15:0] addr_selector3_3342;
wire[15:0] addr_remain3_3342;
address_decode_4 decoder_3_3342 = address_decode_4(addr_selector2_208[14],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3342,addr_remain3_3342);


wire[15:0] addr_selector3_3343;
wire[15:0] addr_remain3_3343;
address_decode_4 decoder_3_3343 = address_decode_4(addr_selector2_208[15],addr_remain2_208[15:0],addr_remain2_208,addr_selector3_3343,addr_remain3_3343);


wire[15:0] addr_selector3_3344;
wire[15:0] addr_remain3_3344;
address_decode_4 decoder_3_3344 = address_decode_4(addr_selector2_209[0],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3344,addr_remain3_3344);


wire[15:0] addr_selector3_3345;
wire[15:0] addr_remain3_3345;
address_decode_4 decoder_3_3345 = address_decode_4(addr_selector2_209[1],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3345,addr_remain3_3345);


wire[15:0] addr_selector3_3346;
wire[15:0] addr_remain3_3346;
address_decode_4 decoder_3_3346 = address_decode_4(addr_selector2_209[2],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3346,addr_remain3_3346);


wire[15:0] addr_selector3_3347;
wire[15:0] addr_remain3_3347;
address_decode_4 decoder_3_3347 = address_decode_4(addr_selector2_209[3],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3347,addr_remain3_3347);


wire[15:0] addr_selector3_3348;
wire[15:0] addr_remain3_3348;
address_decode_4 decoder_3_3348 = address_decode_4(addr_selector2_209[4],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3348,addr_remain3_3348);


wire[15:0] addr_selector3_3349;
wire[15:0] addr_remain3_3349;
address_decode_4 decoder_3_3349 = address_decode_4(addr_selector2_209[5],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3349,addr_remain3_3349);


wire[15:0] addr_selector3_3350;
wire[15:0] addr_remain3_3350;
address_decode_4 decoder_3_3350 = address_decode_4(addr_selector2_209[6],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3350,addr_remain3_3350);


wire[15:0] addr_selector3_3351;
wire[15:0] addr_remain3_3351;
address_decode_4 decoder_3_3351 = address_decode_4(addr_selector2_209[7],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3351,addr_remain3_3351);


wire[15:0] addr_selector3_3352;
wire[15:0] addr_remain3_3352;
address_decode_4 decoder_3_3352 = address_decode_4(addr_selector2_209[8],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3352,addr_remain3_3352);


wire[15:0] addr_selector3_3353;
wire[15:0] addr_remain3_3353;
address_decode_4 decoder_3_3353 = address_decode_4(addr_selector2_209[9],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3353,addr_remain3_3353);


wire[15:0] addr_selector3_3354;
wire[15:0] addr_remain3_3354;
address_decode_4 decoder_3_3354 = address_decode_4(addr_selector2_209[10],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3354,addr_remain3_3354);


wire[15:0] addr_selector3_3355;
wire[15:0] addr_remain3_3355;
address_decode_4 decoder_3_3355 = address_decode_4(addr_selector2_209[11],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3355,addr_remain3_3355);


wire[15:0] addr_selector3_3356;
wire[15:0] addr_remain3_3356;
address_decode_4 decoder_3_3356 = address_decode_4(addr_selector2_209[12],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3356,addr_remain3_3356);


wire[15:0] addr_selector3_3357;
wire[15:0] addr_remain3_3357;
address_decode_4 decoder_3_3357 = address_decode_4(addr_selector2_209[13],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3357,addr_remain3_3357);


wire[15:0] addr_selector3_3358;
wire[15:0] addr_remain3_3358;
address_decode_4 decoder_3_3358 = address_decode_4(addr_selector2_209[14],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3358,addr_remain3_3358);


wire[15:0] addr_selector3_3359;
wire[15:0] addr_remain3_3359;
address_decode_4 decoder_3_3359 = address_decode_4(addr_selector2_209[15],addr_remain2_209[15:0],addr_remain2_209,addr_selector3_3359,addr_remain3_3359);


wire[15:0] addr_selector3_3360;
wire[15:0] addr_remain3_3360;
address_decode_4 decoder_3_3360 = address_decode_4(addr_selector2_210[0],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3360,addr_remain3_3360);


wire[15:0] addr_selector3_3361;
wire[15:0] addr_remain3_3361;
address_decode_4 decoder_3_3361 = address_decode_4(addr_selector2_210[1],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3361,addr_remain3_3361);


wire[15:0] addr_selector3_3362;
wire[15:0] addr_remain3_3362;
address_decode_4 decoder_3_3362 = address_decode_4(addr_selector2_210[2],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3362,addr_remain3_3362);


wire[15:0] addr_selector3_3363;
wire[15:0] addr_remain3_3363;
address_decode_4 decoder_3_3363 = address_decode_4(addr_selector2_210[3],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3363,addr_remain3_3363);


wire[15:0] addr_selector3_3364;
wire[15:0] addr_remain3_3364;
address_decode_4 decoder_3_3364 = address_decode_4(addr_selector2_210[4],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3364,addr_remain3_3364);


wire[15:0] addr_selector3_3365;
wire[15:0] addr_remain3_3365;
address_decode_4 decoder_3_3365 = address_decode_4(addr_selector2_210[5],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3365,addr_remain3_3365);


wire[15:0] addr_selector3_3366;
wire[15:0] addr_remain3_3366;
address_decode_4 decoder_3_3366 = address_decode_4(addr_selector2_210[6],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3366,addr_remain3_3366);


wire[15:0] addr_selector3_3367;
wire[15:0] addr_remain3_3367;
address_decode_4 decoder_3_3367 = address_decode_4(addr_selector2_210[7],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3367,addr_remain3_3367);


wire[15:0] addr_selector3_3368;
wire[15:0] addr_remain3_3368;
address_decode_4 decoder_3_3368 = address_decode_4(addr_selector2_210[8],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3368,addr_remain3_3368);


wire[15:0] addr_selector3_3369;
wire[15:0] addr_remain3_3369;
address_decode_4 decoder_3_3369 = address_decode_4(addr_selector2_210[9],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3369,addr_remain3_3369);


wire[15:0] addr_selector3_3370;
wire[15:0] addr_remain3_3370;
address_decode_4 decoder_3_3370 = address_decode_4(addr_selector2_210[10],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3370,addr_remain3_3370);


wire[15:0] addr_selector3_3371;
wire[15:0] addr_remain3_3371;
address_decode_4 decoder_3_3371 = address_decode_4(addr_selector2_210[11],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3371,addr_remain3_3371);


wire[15:0] addr_selector3_3372;
wire[15:0] addr_remain3_3372;
address_decode_4 decoder_3_3372 = address_decode_4(addr_selector2_210[12],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3372,addr_remain3_3372);


wire[15:0] addr_selector3_3373;
wire[15:0] addr_remain3_3373;
address_decode_4 decoder_3_3373 = address_decode_4(addr_selector2_210[13],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3373,addr_remain3_3373);


wire[15:0] addr_selector3_3374;
wire[15:0] addr_remain3_3374;
address_decode_4 decoder_3_3374 = address_decode_4(addr_selector2_210[14],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3374,addr_remain3_3374);


wire[15:0] addr_selector3_3375;
wire[15:0] addr_remain3_3375;
address_decode_4 decoder_3_3375 = address_decode_4(addr_selector2_210[15],addr_remain2_210[15:0],addr_remain2_210,addr_selector3_3375,addr_remain3_3375);


wire[15:0] addr_selector3_3376;
wire[15:0] addr_remain3_3376;
address_decode_4 decoder_3_3376 = address_decode_4(addr_selector2_211[0],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3376,addr_remain3_3376);


wire[15:0] addr_selector3_3377;
wire[15:0] addr_remain3_3377;
address_decode_4 decoder_3_3377 = address_decode_4(addr_selector2_211[1],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3377,addr_remain3_3377);


wire[15:0] addr_selector3_3378;
wire[15:0] addr_remain3_3378;
address_decode_4 decoder_3_3378 = address_decode_4(addr_selector2_211[2],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3378,addr_remain3_3378);


wire[15:0] addr_selector3_3379;
wire[15:0] addr_remain3_3379;
address_decode_4 decoder_3_3379 = address_decode_4(addr_selector2_211[3],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3379,addr_remain3_3379);


wire[15:0] addr_selector3_3380;
wire[15:0] addr_remain3_3380;
address_decode_4 decoder_3_3380 = address_decode_4(addr_selector2_211[4],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3380,addr_remain3_3380);


wire[15:0] addr_selector3_3381;
wire[15:0] addr_remain3_3381;
address_decode_4 decoder_3_3381 = address_decode_4(addr_selector2_211[5],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3381,addr_remain3_3381);


wire[15:0] addr_selector3_3382;
wire[15:0] addr_remain3_3382;
address_decode_4 decoder_3_3382 = address_decode_4(addr_selector2_211[6],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3382,addr_remain3_3382);


wire[15:0] addr_selector3_3383;
wire[15:0] addr_remain3_3383;
address_decode_4 decoder_3_3383 = address_decode_4(addr_selector2_211[7],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3383,addr_remain3_3383);


wire[15:0] addr_selector3_3384;
wire[15:0] addr_remain3_3384;
address_decode_4 decoder_3_3384 = address_decode_4(addr_selector2_211[8],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3384,addr_remain3_3384);


wire[15:0] addr_selector3_3385;
wire[15:0] addr_remain3_3385;
address_decode_4 decoder_3_3385 = address_decode_4(addr_selector2_211[9],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3385,addr_remain3_3385);


wire[15:0] addr_selector3_3386;
wire[15:0] addr_remain3_3386;
address_decode_4 decoder_3_3386 = address_decode_4(addr_selector2_211[10],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3386,addr_remain3_3386);


wire[15:0] addr_selector3_3387;
wire[15:0] addr_remain3_3387;
address_decode_4 decoder_3_3387 = address_decode_4(addr_selector2_211[11],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3387,addr_remain3_3387);


wire[15:0] addr_selector3_3388;
wire[15:0] addr_remain3_3388;
address_decode_4 decoder_3_3388 = address_decode_4(addr_selector2_211[12],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3388,addr_remain3_3388);


wire[15:0] addr_selector3_3389;
wire[15:0] addr_remain3_3389;
address_decode_4 decoder_3_3389 = address_decode_4(addr_selector2_211[13],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3389,addr_remain3_3389);


wire[15:0] addr_selector3_3390;
wire[15:0] addr_remain3_3390;
address_decode_4 decoder_3_3390 = address_decode_4(addr_selector2_211[14],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3390,addr_remain3_3390);


wire[15:0] addr_selector3_3391;
wire[15:0] addr_remain3_3391;
address_decode_4 decoder_3_3391 = address_decode_4(addr_selector2_211[15],addr_remain2_211[15:0],addr_remain2_211,addr_selector3_3391,addr_remain3_3391);


wire[15:0] addr_selector3_3392;
wire[15:0] addr_remain3_3392;
address_decode_4 decoder_3_3392 = address_decode_4(addr_selector2_212[0],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3392,addr_remain3_3392);


wire[15:0] addr_selector3_3393;
wire[15:0] addr_remain3_3393;
address_decode_4 decoder_3_3393 = address_decode_4(addr_selector2_212[1],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3393,addr_remain3_3393);


wire[15:0] addr_selector3_3394;
wire[15:0] addr_remain3_3394;
address_decode_4 decoder_3_3394 = address_decode_4(addr_selector2_212[2],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3394,addr_remain3_3394);


wire[15:0] addr_selector3_3395;
wire[15:0] addr_remain3_3395;
address_decode_4 decoder_3_3395 = address_decode_4(addr_selector2_212[3],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3395,addr_remain3_3395);


wire[15:0] addr_selector3_3396;
wire[15:0] addr_remain3_3396;
address_decode_4 decoder_3_3396 = address_decode_4(addr_selector2_212[4],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3396,addr_remain3_3396);


wire[15:0] addr_selector3_3397;
wire[15:0] addr_remain3_3397;
address_decode_4 decoder_3_3397 = address_decode_4(addr_selector2_212[5],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3397,addr_remain3_3397);


wire[15:0] addr_selector3_3398;
wire[15:0] addr_remain3_3398;
address_decode_4 decoder_3_3398 = address_decode_4(addr_selector2_212[6],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3398,addr_remain3_3398);


wire[15:0] addr_selector3_3399;
wire[15:0] addr_remain3_3399;
address_decode_4 decoder_3_3399 = address_decode_4(addr_selector2_212[7],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3399,addr_remain3_3399);


wire[15:0] addr_selector3_3400;
wire[15:0] addr_remain3_3400;
address_decode_4 decoder_3_3400 = address_decode_4(addr_selector2_212[8],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3400,addr_remain3_3400);


wire[15:0] addr_selector3_3401;
wire[15:0] addr_remain3_3401;
address_decode_4 decoder_3_3401 = address_decode_4(addr_selector2_212[9],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3401,addr_remain3_3401);


wire[15:0] addr_selector3_3402;
wire[15:0] addr_remain3_3402;
address_decode_4 decoder_3_3402 = address_decode_4(addr_selector2_212[10],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3402,addr_remain3_3402);


wire[15:0] addr_selector3_3403;
wire[15:0] addr_remain3_3403;
address_decode_4 decoder_3_3403 = address_decode_4(addr_selector2_212[11],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3403,addr_remain3_3403);


wire[15:0] addr_selector3_3404;
wire[15:0] addr_remain3_3404;
address_decode_4 decoder_3_3404 = address_decode_4(addr_selector2_212[12],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3404,addr_remain3_3404);


wire[15:0] addr_selector3_3405;
wire[15:0] addr_remain3_3405;
address_decode_4 decoder_3_3405 = address_decode_4(addr_selector2_212[13],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3405,addr_remain3_3405);


wire[15:0] addr_selector3_3406;
wire[15:0] addr_remain3_3406;
address_decode_4 decoder_3_3406 = address_decode_4(addr_selector2_212[14],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3406,addr_remain3_3406);


wire[15:0] addr_selector3_3407;
wire[15:0] addr_remain3_3407;
address_decode_4 decoder_3_3407 = address_decode_4(addr_selector2_212[15],addr_remain2_212[15:0],addr_remain2_212,addr_selector3_3407,addr_remain3_3407);


wire[15:0] addr_selector3_3408;
wire[15:0] addr_remain3_3408;
address_decode_4 decoder_3_3408 = address_decode_4(addr_selector2_213[0],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3408,addr_remain3_3408);


wire[15:0] addr_selector3_3409;
wire[15:0] addr_remain3_3409;
address_decode_4 decoder_3_3409 = address_decode_4(addr_selector2_213[1],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3409,addr_remain3_3409);


wire[15:0] addr_selector3_3410;
wire[15:0] addr_remain3_3410;
address_decode_4 decoder_3_3410 = address_decode_4(addr_selector2_213[2],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3410,addr_remain3_3410);


wire[15:0] addr_selector3_3411;
wire[15:0] addr_remain3_3411;
address_decode_4 decoder_3_3411 = address_decode_4(addr_selector2_213[3],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3411,addr_remain3_3411);


wire[15:0] addr_selector3_3412;
wire[15:0] addr_remain3_3412;
address_decode_4 decoder_3_3412 = address_decode_4(addr_selector2_213[4],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3412,addr_remain3_3412);


wire[15:0] addr_selector3_3413;
wire[15:0] addr_remain3_3413;
address_decode_4 decoder_3_3413 = address_decode_4(addr_selector2_213[5],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3413,addr_remain3_3413);


wire[15:0] addr_selector3_3414;
wire[15:0] addr_remain3_3414;
address_decode_4 decoder_3_3414 = address_decode_4(addr_selector2_213[6],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3414,addr_remain3_3414);


wire[15:0] addr_selector3_3415;
wire[15:0] addr_remain3_3415;
address_decode_4 decoder_3_3415 = address_decode_4(addr_selector2_213[7],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3415,addr_remain3_3415);


wire[15:0] addr_selector3_3416;
wire[15:0] addr_remain3_3416;
address_decode_4 decoder_3_3416 = address_decode_4(addr_selector2_213[8],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3416,addr_remain3_3416);


wire[15:0] addr_selector3_3417;
wire[15:0] addr_remain3_3417;
address_decode_4 decoder_3_3417 = address_decode_4(addr_selector2_213[9],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3417,addr_remain3_3417);


wire[15:0] addr_selector3_3418;
wire[15:0] addr_remain3_3418;
address_decode_4 decoder_3_3418 = address_decode_4(addr_selector2_213[10],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3418,addr_remain3_3418);


wire[15:0] addr_selector3_3419;
wire[15:0] addr_remain3_3419;
address_decode_4 decoder_3_3419 = address_decode_4(addr_selector2_213[11],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3419,addr_remain3_3419);


wire[15:0] addr_selector3_3420;
wire[15:0] addr_remain3_3420;
address_decode_4 decoder_3_3420 = address_decode_4(addr_selector2_213[12],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3420,addr_remain3_3420);


wire[15:0] addr_selector3_3421;
wire[15:0] addr_remain3_3421;
address_decode_4 decoder_3_3421 = address_decode_4(addr_selector2_213[13],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3421,addr_remain3_3421);


wire[15:0] addr_selector3_3422;
wire[15:0] addr_remain3_3422;
address_decode_4 decoder_3_3422 = address_decode_4(addr_selector2_213[14],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3422,addr_remain3_3422);


wire[15:0] addr_selector3_3423;
wire[15:0] addr_remain3_3423;
address_decode_4 decoder_3_3423 = address_decode_4(addr_selector2_213[15],addr_remain2_213[15:0],addr_remain2_213,addr_selector3_3423,addr_remain3_3423);


wire[15:0] addr_selector3_3424;
wire[15:0] addr_remain3_3424;
address_decode_4 decoder_3_3424 = address_decode_4(addr_selector2_214[0],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3424,addr_remain3_3424);


wire[15:0] addr_selector3_3425;
wire[15:0] addr_remain3_3425;
address_decode_4 decoder_3_3425 = address_decode_4(addr_selector2_214[1],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3425,addr_remain3_3425);


wire[15:0] addr_selector3_3426;
wire[15:0] addr_remain3_3426;
address_decode_4 decoder_3_3426 = address_decode_4(addr_selector2_214[2],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3426,addr_remain3_3426);


wire[15:0] addr_selector3_3427;
wire[15:0] addr_remain3_3427;
address_decode_4 decoder_3_3427 = address_decode_4(addr_selector2_214[3],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3427,addr_remain3_3427);


wire[15:0] addr_selector3_3428;
wire[15:0] addr_remain3_3428;
address_decode_4 decoder_3_3428 = address_decode_4(addr_selector2_214[4],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3428,addr_remain3_3428);


wire[15:0] addr_selector3_3429;
wire[15:0] addr_remain3_3429;
address_decode_4 decoder_3_3429 = address_decode_4(addr_selector2_214[5],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3429,addr_remain3_3429);


wire[15:0] addr_selector3_3430;
wire[15:0] addr_remain3_3430;
address_decode_4 decoder_3_3430 = address_decode_4(addr_selector2_214[6],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3430,addr_remain3_3430);


wire[15:0] addr_selector3_3431;
wire[15:0] addr_remain3_3431;
address_decode_4 decoder_3_3431 = address_decode_4(addr_selector2_214[7],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3431,addr_remain3_3431);


wire[15:0] addr_selector3_3432;
wire[15:0] addr_remain3_3432;
address_decode_4 decoder_3_3432 = address_decode_4(addr_selector2_214[8],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3432,addr_remain3_3432);


wire[15:0] addr_selector3_3433;
wire[15:0] addr_remain3_3433;
address_decode_4 decoder_3_3433 = address_decode_4(addr_selector2_214[9],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3433,addr_remain3_3433);


wire[15:0] addr_selector3_3434;
wire[15:0] addr_remain3_3434;
address_decode_4 decoder_3_3434 = address_decode_4(addr_selector2_214[10],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3434,addr_remain3_3434);


wire[15:0] addr_selector3_3435;
wire[15:0] addr_remain3_3435;
address_decode_4 decoder_3_3435 = address_decode_4(addr_selector2_214[11],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3435,addr_remain3_3435);


wire[15:0] addr_selector3_3436;
wire[15:0] addr_remain3_3436;
address_decode_4 decoder_3_3436 = address_decode_4(addr_selector2_214[12],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3436,addr_remain3_3436);


wire[15:0] addr_selector3_3437;
wire[15:0] addr_remain3_3437;
address_decode_4 decoder_3_3437 = address_decode_4(addr_selector2_214[13],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3437,addr_remain3_3437);


wire[15:0] addr_selector3_3438;
wire[15:0] addr_remain3_3438;
address_decode_4 decoder_3_3438 = address_decode_4(addr_selector2_214[14],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3438,addr_remain3_3438);


wire[15:0] addr_selector3_3439;
wire[15:0] addr_remain3_3439;
address_decode_4 decoder_3_3439 = address_decode_4(addr_selector2_214[15],addr_remain2_214[15:0],addr_remain2_214,addr_selector3_3439,addr_remain3_3439);


wire[15:0] addr_selector3_3440;
wire[15:0] addr_remain3_3440;
address_decode_4 decoder_3_3440 = address_decode_4(addr_selector2_215[0],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3440,addr_remain3_3440);


wire[15:0] addr_selector3_3441;
wire[15:0] addr_remain3_3441;
address_decode_4 decoder_3_3441 = address_decode_4(addr_selector2_215[1],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3441,addr_remain3_3441);


wire[15:0] addr_selector3_3442;
wire[15:0] addr_remain3_3442;
address_decode_4 decoder_3_3442 = address_decode_4(addr_selector2_215[2],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3442,addr_remain3_3442);


wire[15:0] addr_selector3_3443;
wire[15:0] addr_remain3_3443;
address_decode_4 decoder_3_3443 = address_decode_4(addr_selector2_215[3],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3443,addr_remain3_3443);


wire[15:0] addr_selector3_3444;
wire[15:0] addr_remain3_3444;
address_decode_4 decoder_3_3444 = address_decode_4(addr_selector2_215[4],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3444,addr_remain3_3444);


wire[15:0] addr_selector3_3445;
wire[15:0] addr_remain3_3445;
address_decode_4 decoder_3_3445 = address_decode_4(addr_selector2_215[5],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3445,addr_remain3_3445);


wire[15:0] addr_selector3_3446;
wire[15:0] addr_remain3_3446;
address_decode_4 decoder_3_3446 = address_decode_4(addr_selector2_215[6],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3446,addr_remain3_3446);


wire[15:0] addr_selector3_3447;
wire[15:0] addr_remain3_3447;
address_decode_4 decoder_3_3447 = address_decode_4(addr_selector2_215[7],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3447,addr_remain3_3447);


wire[15:0] addr_selector3_3448;
wire[15:0] addr_remain3_3448;
address_decode_4 decoder_3_3448 = address_decode_4(addr_selector2_215[8],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3448,addr_remain3_3448);


wire[15:0] addr_selector3_3449;
wire[15:0] addr_remain3_3449;
address_decode_4 decoder_3_3449 = address_decode_4(addr_selector2_215[9],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3449,addr_remain3_3449);


wire[15:0] addr_selector3_3450;
wire[15:0] addr_remain3_3450;
address_decode_4 decoder_3_3450 = address_decode_4(addr_selector2_215[10],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3450,addr_remain3_3450);


wire[15:0] addr_selector3_3451;
wire[15:0] addr_remain3_3451;
address_decode_4 decoder_3_3451 = address_decode_4(addr_selector2_215[11],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3451,addr_remain3_3451);


wire[15:0] addr_selector3_3452;
wire[15:0] addr_remain3_3452;
address_decode_4 decoder_3_3452 = address_decode_4(addr_selector2_215[12],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3452,addr_remain3_3452);


wire[15:0] addr_selector3_3453;
wire[15:0] addr_remain3_3453;
address_decode_4 decoder_3_3453 = address_decode_4(addr_selector2_215[13],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3453,addr_remain3_3453);


wire[15:0] addr_selector3_3454;
wire[15:0] addr_remain3_3454;
address_decode_4 decoder_3_3454 = address_decode_4(addr_selector2_215[14],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3454,addr_remain3_3454);


wire[15:0] addr_selector3_3455;
wire[15:0] addr_remain3_3455;
address_decode_4 decoder_3_3455 = address_decode_4(addr_selector2_215[15],addr_remain2_215[15:0],addr_remain2_215,addr_selector3_3455,addr_remain3_3455);


wire[15:0] addr_selector3_3456;
wire[15:0] addr_remain3_3456;
address_decode_4 decoder_3_3456 = address_decode_4(addr_selector2_216[0],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3456,addr_remain3_3456);


wire[15:0] addr_selector3_3457;
wire[15:0] addr_remain3_3457;
address_decode_4 decoder_3_3457 = address_decode_4(addr_selector2_216[1],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3457,addr_remain3_3457);


wire[15:0] addr_selector3_3458;
wire[15:0] addr_remain3_3458;
address_decode_4 decoder_3_3458 = address_decode_4(addr_selector2_216[2],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3458,addr_remain3_3458);


wire[15:0] addr_selector3_3459;
wire[15:0] addr_remain3_3459;
address_decode_4 decoder_3_3459 = address_decode_4(addr_selector2_216[3],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3459,addr_remain3_3459);


wire[15:0] addr_selector3_3460;
wire[15:0] addr_remain3_3460;
address_decode_4 decoder_3_3460 = address_decode_4(addr_selector2_216[4],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3460,addr_remain3_3460);


wire[15:0] addr_selector3_3461;
wire[15:0] addr_remain3_3461;
address_decode_4 decoder_3_3461 = address_decode_4(addr_selector2_216[5],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3461,addr_remain3_3461);


wire[15:0] addr_selector3_3462;
wire[15:0] addr_remain3_3462;
address_decode_4 decoder_3_3462 = address_decode_4(addr_selector2_216[6],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3462,addr_remain3_3462);


wire[15:0] addr_selector3_3463;
wire[15:0] addr_remain3_3463;
address_decode_4 decoder_3_3463 = address_decode_4(addr_selector2_216[7],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3463,addr_remain3_3463);


wire[15:0] addr_selector3_3464;
wire[15:0] addr_remain3_3464;
address_decode_4 decoder_3_3464 = address_decode_4(addr_selector2_216[8],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3464,addr_remain3_3464);


wire[15:0] addr_selector3_3465;
wire[15:0] addr_remain3_3465;
address_decode_4 decoder_3_3465 = address_decode_4(addr_selector2_216[9],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3465,addr_remain3_3465);


wire[15:0] addr_selector3_3466;
wire[15:0] addr_remain3_3466;
address_decode_4 decoder_3_3466 = address_decode_4(addr_selector2_216[10],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3466,addr_remain3_3466);


wire[15:0] addr_selector3_3467;
wire[15:0] addr_remain3_3467;
address_decode_4 decoder_3_3467 = address_decode_4(addr_selector2_216[11],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3467,addr_remain3_3467);


wire[15:0] addr_selector3_3468;
wire[15:0] addr_remain3_3468;
address_decode_4 decoder_3_3468 = address_decode_4(addr_selector2_216[12],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3468,addr_remain3_3468);


wire[15:0] addr_selector3_3469;
wire[15:0] addr_remain3_3469;
address_decode_4 decoder_3_3469 = address_decode_4(addr_selector2_216[13],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3469,addr_remain3_3469);


wire[15:0] addr_selector3_3470;
wire[15:0] addr_remain3_3470;
address_decode_4 decoder_3_3470 = address_decode_4(addr_selector2_216[14],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3470,addr_remain3_3470);


wire[15:0] addr_selector3_3471;
wire[15:0] addr_remain3_3471;
address_decode_4 decoder_3_3471 = address_decode_4(addr_selector2_216[15],addr_remain2_216[15:0],addr_remain2_216,addr_selector3_3471,addr_remain3_3471);


wire[15:0] addr_selector3_3472;
wire[15:0] addr_remain3_3472;
address_decode_4 decoder_3_3472 = address_decode_4(addr_selector2_217[0],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3472,addr_remain3_3472);


wire[15:0] addr_selector3_3473;
wire[15:0] addr_remain3_3473;
address_decode_4 decoder_3_3473 = address_decode_4(addr_selector2_217[1],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3473,addr_remain3_3473);


wire[15:0] addr_selector3_3474;
wire[15:0] addr_remain3_3474;
address_decode_4 decoder_3_3474 = address_decode_4(addr_selector2_217[2],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3474,addr_remain3_3474);


wire[15:0] addr_selector3_3475;
wire[15:0] addr_remain3_3475;
address_decode_4 decoder_3_3475 = address_decode_4(addr_selector2_217[3],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3475,addr_remain3_3475);


wire[15:0] addr_selector3_3476;
wire[15:0] addr_remain3_3476;
address_decode_4 decoder_3_3476 = address_decode_4(addr_selector2_217[4],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3476,addr_remain3_3476);


wire[15:0] addr_selector3_3477;
wire[15:0] addr_remain3_3477;
address_decode_4 decoder_3_3477 = address_decode_4(addr_selector2_217[5],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3477,addr_remain3_3477);


wire[15:0] addr_selector3_3478;
wire[15:0] addr_remain3_3478;
address_decode_4 decoder_3_3478 = address_decode_4(addr_selector2_217[6],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3478,addr_remain3_3478);


wire[15:0] addr_selector3_3479;
wire[15:0] addr_remain3_3479;
address_decode_4 decoder_3_3479 = address_decode_4(addr_selector2_217[7],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3479,addr_remain3_3479);


wire[15:0] addr_selector3_3480;
wire[15:0] addr_remain3_3480;
address_decode_4 decoder_3_3480 = address_decode_4(addr_selector2_217[8],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3480,addr_remain3_3480);


wire[15:0] addr_selector3_3481;
wire[15:0] addr_remain3_3481;
address_decode_4 decoder_3_3481 = address_decode_4(addr_selector2_217[9],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3481,addr_remain3_3481);


wire[15:0] addr_selector3_3482;
wire[15:0] addr_remain3_3482;
address_decode_4 decoder_3_3482 = address_decode_4(addr_selector2_217[10],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3482,addr_remain3_3482);


wire[15:0] addr_selector3_3483;
wire[15:0] addr_remain3_3483;
address_decode_4 decoder_3_3483 = address_decode_4(addr_selector2_217[11],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3483,addr_remain3_3483);


wire[15:0] addr_selector3_3484;
wire[15:0] addr_remain3_3484;
address_decode_4 decoder_3_3484 = address_decode_4(addr_selector2_217[12],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3484,addr_remain3_3484);


wire[15:0] addr_selector3_3485;
wire[15:0] addr_remain3_3485;
address_decode_4 decoder_3_3485 = address_decode_4(addr_selector2_217[13],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3485,addr_remain3_3485);


wire[15:0] addr_selector3_3486;
wire[15:0] addr_remain3_3486;
address_decode_4 decoder_3_3486 = address_decode_4(addr_selector2_217[14],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3486,addr_remain3_3486);


wire[15:0] addr_selector3_3487;
wire[15:0] addr_remain3_3487;
address_decode_4 decoder_3_3487 = address_decode_4(addr_selector2_217[15],addr_remain2_217[15:0],addr_remain2_217,addr_selector3_3487,addr_remain3_3487);


wire[15:0] addr_selector3_3488;
wire[15:0] addr_remain3_3488;
address_decode_4 decoder_3_3488 = address_decode_4(addr_selector2_218[0],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3488,addr_remain3_3488);


wire[15:0] addr_selector3_3489;
wire[15:0] addr_remain3_3489;
address_decode_4 decoder_3_3489 = address_decode_4(addr_selector2_218[1],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3489,addr_remain3_3489);


wire[15:0] addr_selector3_3490;
wire[15:0] addr_remain3_3490;
address_decode_4 decoder_3_3490 = address_decode_4(addr_selector2_218[2],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3490,addr_remain3_3490);


wire[15:0] addr_selector3_3491;
wire[15:0] addr_remain3_3491;
address_decode_4 decoder_3_3491 = address_decode_4(addr_selector2_218[3],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3491,addr_remain3_3491);


wire[15:0] addr_selector3_3492;
wire[15:0] addr_remain3_3492;
address_decode_4 decoder_3_3492 = address_decode_4(addr_selector2_218[4],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3492,addr_remain3_3492);


wire[15:0] addr_selector3_3493;
wire[15:0] addr_remain3_3493;
address_decode_4 decoder_3_3493 = address_decode_4(addr_selector2_218[5],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3493,addr_remain3_3493);


wire[15:0] addr_selector3_3494;
wire[15:0] addr_remain3_3494;
address_decode_4 decoder_3_3494 = address_decode_4(addr_selector2_218[6],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3494,addr_remain3_3494);


wire[15:0] addr_selector3_3495;
wire[15:0] addr_remain3_3495;
address_decode_4 decoder_3_3495 = address_decode_4(addr_selector2_218[7],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3495,addr_remain3_3495);


wire[15:0] addr_selector3_3496;
wire[15:0] addr_remain3_3496;
address_decode_4 decoder_3_3496 = address_decode_4(addr_selector2_218[8],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3496,addr_remain3_3496);


wire[15:0] addr_selector3_3497;
wire[15:0] addr_remain3_3497;
address_decode_4 decoder_3_3497 = address_decode_4(addr_selector2_218[9],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3497,addr_remain3_3497);


wire[15:0] addr_selector3_3498;
wire[15:0] addr_remain3_3498;
address_decode_4 decoder_3_3498 = address_decode_4(addr_selector2_218[10],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3498,addr_remain3_3498);


wire[15:0] addr_selector3_3499;
wire[15:0] addr_remain3_3499;
address_decode_4 decoder_3_3499 = address_decode_4(addr_selector2_218[11],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3499,addr_remain3_3499);


wire[15:0] addr_selector3_3500;
wire[15:0] addr_remain3_3500;
address_decode_4 decoder_3_3500 = address_decode_4(addr_selector2_218[12],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3500,addr_remain3_3500);


wire[15:0] addr_selector3_3501;
wire[15:0] addr_remain3_3501;
address_decode_4 decoder_3_3501 = address_decode_4(addr_selector2_218[13],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3501,addr_remain3_3501);


wire[15:0] addr_selector3_3502;
wire[15:0] addr_remain3_3502;
address_decode_4 decoder_3_3502 = address_decode_4(addr_selector2_218[14],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3502,addr_remain3_3502);


wire[15:0] addr_selector3_3503;
wire[15:0] addr_remain3_3503;
address_decode_4 decoder_3_3503 = address_decode_4(addr_selector2_218[15],addr_remain2_218[15:0],addr_remain2_218,addr_selector3_3503,addr_remain3_3503);


wire[15:0] addr_selector3_3504;
wire[15:0] addr_remain3_3504;
address_decode_4 decoder_3_3504 = address_decode_4(addr_selector2_219[0],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3504,addr_remain3_3504);


wire[15:0] addr_selector3_3505;
wire[15:0] addr_remain3_3505;
address_decode_4 decoder_3_3505 = address_decode_4(addr_selector2_219[1],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3505,addr_remain3_3505);


wire[15:0] addr_selector3_3506;
wire[15:0] addr_remain3_3506;
address_decode_4 decoder_3_3506 = address_decode_4(addr_selector2_219[2],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3506,addr_remain3_3506);


wire[15:0] addr_selector3_3507;
wire[15:0] addr_remain3_3507;
address_decode_4 decoder_3_3507 = address_decode_4(addr_selector2_219[3],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3507,addr_remain3_3507);


wire[15:0] addr_selector3_3508;
wire[15:0] addr_remain3_3508;
address_decode_4 decoder_3_3508 = address_decode_4(addr_selector2_219[4],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3508,addr_remain3_3508);


wire[15:0] addr_selector3_3509;
wire[15:0] addr_remain3_3509;
address_decode_4 decoder_3_3509 = address_decode_4(addr_selector2_219[5],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3509,addr_remain3_3509);


wire[15:0] addr_selector3_3510;
wire[15:0] addr_remain3_3510;
address_decode_4 decoder_3_3510 = address_decode_4(addr_selector2_219[6],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3510,addr_remain3_3510);


wire[15:0] addr_selector3_3511;
wire[15:0] addr_remain3_3511;
address_decode_4 decoder_3_3511 = address_decode_4(addr_selector2_219[7],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3511,addr_remain3_3511);


wire[15:0] addr_selector3_3512;
wire[15:0] addr_remain3_3512;
address_decode_4 decoder_3_3512 = address_decode_4(addr_selector2_219[8],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3512,addr_remain3_3512);


wire[15:0] addr_selector3_3513;
wire[15:0] addr_remain3_3513;
address_decode_4 decoder_3_3513 = address_decode_4(addr_selector2_219[9],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3513,addr_remain3_3513);


wire[15:0] addr_selector3_3514;
wire[15:0] addr_remain3_3514;
address_decode_4 decoder_3_3514 = address_decode_4(addr_selector2_219[10],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3514,addr_remain3_3514);


wire[15:0] addr_selector3_3515;
wire[15:0] addr_remain3_3515;
address_decode_4 decoder_3_3515 = address_decode_4(addr_selector2_219[11],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3515,addr_remain3_3515);


wire[15:0] addr_selector3_3516;
wire[15:0] addr_remain3_3516;
address_decode_4 decoder_3_3516 = address_decode_4(addr_selector2_219[12],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3516,addr_remain3_3516);


wire[15:0] addr_selector3_3517;
wire[15:0] addr_remain3_3517;
address_decode_4 decoder_3_3517 = address_decode_4(addr_selector2_219[13],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3517,addr_remain3_3517);


wire[15:0] addr_selector3_3518;
wire[15:0] addr_remain3_3518;
address_decode_4 decoder_3_3518 = address_decode_4(addr_selector2_219[14],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3518,addr_remain3_3518);


wire[15:0] addr_selector3_3519;
wire[15:0] addr_remain3_3519;
address_decode_4 decoder_3_3519 = address_decode_4(addr_selector2_219[15],addr_remain2_219[15:0],addr_remain2_219,addr_selector3_3519,addr_remain3_3519);


wire[15:0] addr_selector3_3520;
wire[15:0] addr_remain3_3520;
address_decode_4 decoder_3_3520 = address_decode_4(addr_selector2_220[0],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3520,addr_remain3_3520);


wire[15:0] addr_selector3_3521;
wire[15:0] addr_remain3_3521;
address_decode_4 decoder_3_3521 = address_decode_4(addr_selector2_220[1],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3521,addr_remain3_3521);


wire[15:0] addr_selector3_3522;
wire[15:0] addr_remain3_3522;
address_decode_4 decoder_3_3522 = address_decode_4(addr_selector2_220[2],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3522,addr_remain3_3522);


wire[15:0] addr_selector3_3523;
wire[15:0] addr_remain3_3523;
address_decode_4 decoder_3_3523 = address_decode_4(addr_selector2_220[3],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3523,addr_remain3_3523);


wire[15:0] addr_selector3_3524;
wire[15:0] addr_remain3_3524;
address_decode_4 decoder_3_3524 = address_decode_4(addr_selector2_220[4],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3524,addr_remain3_3524);


wire[15:0] addr_selector3_3525;
wire[15:0] addr_remain3_3525;
address_decode_4 decoder_3_3525 = address_decode_4(addr_selector2_220[5],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3525,addr_remain3_3525);


wire[15:0] addr_selector3_3526;
wire[15:0] addr_remain3_3526;
address_decode_4 decoder_3_3526 = address_decode_4(addr_selector2_220[6],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3526,addr_remain3_3526);


wire[15:0] addr_selector3_3527;
wire[15:0] addr_remain3_3527;
address_decode_4 decoder_3_3527 = address_decode_4(addr_selector2_220[7],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3527,addr_remain3_3527);


wire[15:0] addr_selector3_3528;
wire[15:0] addr_remain3_3528;
address_decode_4 decoder_3_3528 = address_decode_4(addr_selector2_220[8],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3528,addr_remain3_3528);


wire[15:0] addr_selector3_3529;
wire[15:0] addr_remain3_3529;
address_decode_4 decoder_3_3529 = address_decode_4(addr_selector2_220[9],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3529,addr_remain3_3529);


wire[15:0] addr_selector3_3530;
wire[15:0] addr_remain3_3530;
address_decode_4 decoder_3_3530 = address_decode_4(addr_selector2_220[10],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3530,addr_remain3_3530);


wire[15:0] addr_selector3_3531;
wire[15:0] addr_remain3_3531;
address_decode_4 decoder_3_3531 = address_decode_4(addr_selector2_220[11],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3531,addr_remain3_3531);


wire[15:0] addr_selector3_3532;
wire[15:0] addr_remain3_3532;
address_decode_4 decoder_3_3532 = address_decode_4(addr_selector2_220[12],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3532,addr_remain3_3532);


wire[15:0] addr_selector3_3533;
wire[15:0] addr_remain3_3533;
address_decode_4 decoder_3_3533 = address_decode_4(addr_selector2_220[13],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3533,addr_remain3_3533);


wire[15:0] addr_selector3_3534;
wire[15:0] addr_remain3_3534;
address_decode_4 decoder_3_3534 = address_decode_4(addr_selector2_220[14],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3534,addr_remain3_3534);


wire[15:0] addr_selector3_3535;
wire[15:0] addr_remain3_3535;
address_decode_4 decoder_3_3535 = address_decode_4(addr_selector2_220[15],addr_remain2_220[15:0],addr_remain2_220,addr_selector3_3535,addr_remain3_3535);


wire[15:0] addr_selector3_3536;
wire[15:0] addr_remain3_3536;
address_decode_4 decoder_3_3536 = address_decode_4(addr_selector2_221[0],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3536,addr_remain3_3536);


wire[15:0] addr_selector3_3537;
wire[15:0] addr_remain3_3537;
address_decode_4 decoder_3_3537 = address_decode_4(addr_selector2_221[1],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3537,addr_remain3_3537);


wire[15:0] addr_selector3_3538;
wire[15:0] addr_remain3_3538;
address_decode_4 decoder_3_3538 = address_decode_4(addr_selector2_221[2],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3538,addr_remain3_3538);


wire[15:0] addr_selector3_3539;
wire[15:0] addr_remain3_3539;
address_decode_4 decoder_3_3539 = address_decode_4(addr_selector2_221[3],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3539,addr_remain3_3539);


wire[15:0] addr_selector3_3540;
wire[15:0] addr_remain3_3540;
address_decode_4 decoder_3_3540 = address_decode_4(addr_selector2_221[4],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3540,addr_remain3_3540);


wire[15:0] addr_selector3_3541;
wire[15:0] addr_remain3_3541;
address_decode_4 decoder_3_3541 = address_decode_4(addr_selector2_221[5],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3541,addr_remain3_3541);


wire[15:0] addr_selector3_3542;
wire[15:0] addr_remain3_3542;
address_decode_4 decoder_3_3542 = address_decode_4(addr_selector2_221[6],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3542,addr_remain3_3542);


wire[15:0] addr_selector3_3543;
wire[15:0] addr_remain3_3543;
address_decode_4 decoder_3_3543 = address_decode_4(addr_selector2_221[7],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3543,addr_remain3_3543);


wire[15:0] addr_selector3_3544;
wire[15:0] addr_remain3_3544;
address_decode_4 decoder_3_3544 = address_decode_4(addr_selector2_221[8],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3544,addr_remain3_3544);


wire[15:0] addr_selector3_3545;
wire[15:0] addr_remain3_3545;
address_decode_4 decoder_3_3545 = address_decode_4(addr_selector2_221[9],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3545,addr_remain3_3545);


wire[15:0] addr_selector3_3546;
wire[15:0] addr_remain3_3546;
address_decode_4 decoder_3_3546 = address_decode_4(addr_selector2_221[10],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3546,addr_remain3_3546);


wire[15:0] addr_selector3_3547;
wire[15:0] addr_remain3_3547;
address_decode_4 decoder_3_3547 = address_decode_4(addr_selector2_221[11],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3547,addr_remain3_3547);


wire[15:0] addr_selector3_3548;
wire[15:0] addr_remain3_3548;
address_decode_4 decoder_3_3548 = address_decode_4(addr_selector2_221[12],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3548,addr_remain3_3548);


wire[15:0] addr_selector3_3549;
wire[15:0] addr_remain3_3549;
address_decode_4 decoder_3_3549 = address_decode_4(addr_selector2_221[13],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3549,addr_remain3_3549);


wire[15:0] addr_selector3_3550;
wire[15:0] addr_remain3_3550;
address_decode_4 decoder_3_3550 = address_decode_4(addr_selector2_221[14],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3550,addr_remain3_3550);


wire[15:0] addr_selector3_3551;
wire[15:0] addr_remain3_3551;
address_decode_4 decoder_3_3551 = address_decode_4(addr_selector2_221[15],addr_remain2_221[15:0],addr_remain2_221,addr_selector3_3551,addr_remain3_3551);


wire[15:0] addr_selector3_3552;
wire[15:0] addr_remain3_3552;
address_decode_4 decoder_3_3552 = address_decode_4(addr_selector2_222[0],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3552,addr_remain3_3552);


wire[15:0] addr_selector3_3553;
wire[15:0] addr_remain3_3553;
address_decode_4 decoder_3_3553 = address_decode_4(addr_selector2_222[1],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3553,addr_remain3_3553);


wire[15:0] addr_selector3_3554;
wire[15:0] addr_remain3_3554;
address_decode_4 decoder_3_3554 = address_decode_4(addr_selector2_222[2],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3554,addr_remain3_3554);


wire[15:0] addr_selector3_3555;
wire[15:0] addr_remain3_3555;
address_decode_4 decoder_3_3555 = address_decode_4(addr_selector2_222[3],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3555,addr_remain3_3555);


wire[15:0] addr_selector3_3556;
wire[15:0] addr_remain3_3556;
address_decode_4 decoder_3_3556 = address_decode_4(addr_selector2_222[4],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3556,addr_remain3_3556);


wire[15:0] addr_selector3_3557;
wire[15:0] addr_remain3_3557;
address_decode_4 decoder_3_3557 = address_decode_4(addr_selector2_222[5],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3557,addr_remain3_3557);


wire[15:0] addr_selector3_3558;
wire[15:0] addr_remain3_3558;
address_decode_4 decoder_3_3558 = address_decode_4(addr_selector2_222[6],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3558,addr_remain3_3558);


wire[15:0] addr_selector3_3559;
wire[15:0] addr_remain3_3559;
address_decode_4 decoder_3_3559 = address_decode_4(addr_selector2_222[7],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3559,addr_remain3_3559);


wire[15:0] addr_selector3_3560;
wire[15:0] addr_remain3_3560;
address_decode_4 decoder_3_3560 = address_decode_4(addr_selector2_222[8],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3560,addr_remain3_3560);


wire[15:0] addr_selector3_3561;
wire[15:0] addr_remain3_3561;
address_decode_4 decoder_3_3561 = address_decode_4(addr_selector2_222[9],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3561,addr_remain3_3561);


wire[15:0] addr_selector3_3562;
wire[15:0] addr_remain3_3562;
address_decode_4 decoder_3_3562 = address_decode_4(addr_selector2_222[10],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3562,addr_remain3_3562);


wire[15:0] addr_selector3_3563;
wire[15:0] addr_remain3_3563;
address_decode_4 decoder_3_3563 = address_decode_4(addr_selector2_222[11],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3563,addr_remain3_3563);


wire[15:0] addr_selector3_3564;
wire[15:0] addr_remain3_3564;
address_decode_4 decoder_3_3564 = address_decode_4(addr_selector2_222[12],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3564,addr_remain3_3564);


wire[15:0] addr_selector3_3565;
wire[15:0] addr_remain3_3565;
address_decode_4 decoder_3_3565 = address_decode_4(addr_selector2_222[13],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3565,addr_remain3_3565);


wire[15:0] addr_selector3_3566;
wire[15:0] addr_remain3_3566;
address_decode_4 decoder_3_3566 = address_decode_4(addr_selector2_222[14],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3566,addr_remain3_3566);


wire[15:0] addr_selector3_3567;
wire[15:0] addr_remain3_3567;
address_decode_4 decoder_3_3567 = address_decode_4(addr_selector2_222[15],addr_remain2_222[15:0],addr_remain2_222,addr_selector3_3567,addr_remain3_3567);


wire[15:0] addr_selector3_3568;
wire[15:0] addr_remain3_3568;
address_decode_4 decoder_3_3568 = address_decode_4(addr_selector2_223[0],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3568,addr_remain3_3568);


wire[15:0] addr_selector3_3569;
wire[15:0] addr_remain3_3569;
address_decode_4 decoder_3_3569 = address_decode_4(addr_selector2_223[1],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3569,addr_remain3_3569);


wire[15:0] addr_selector3_3570;
wire[15:0] addr_remain3_3570;
address_decode_4 decoder_3_3570 = address_decode_4(addr_selector2_223[2],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3570,addr_remain3_3570);


wire[15:0] addr_selector3_3571;
wire[15:0] addr_remain3_3571;
address_decode_4 decoder_3_3571 = address_decode_4(addr_selector2_223[3],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3571,addr_remain3_3571);


wire[15:0] addr_selector3_3572;
wire[15:0] addr_remain3_3572;
address_decode_4 decoder_3_3572 = address_decode_4(addr_selector2_223[4],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3572,addr_remain3_3572);


wire[15:0] addr_selector3_3573;
wire[15:0] addr_remain3_3573;
address_decode_4 decoder_3_3573 = address_decode_4(addr_selector2_223[5],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3573,addr_remain3_3573);


wire[15:0] addr_selector3_3574;
wire[15:0] addr_remain3_3574;
address_decode_4 decoder_3_3574 = address_decode_4(addr_selector2_223[6],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3574,addr_remain3_3574);


wire[15:0] addr_selector3_3575;
wire[15:0] addr_remain3_3575;
address_decode_4 decoder_3_3575 = address_decode_4(addr_selector2_223[7],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3575,addr_remain3_3575);


wire[15:0] addr_selector3_3576;
wire[15:0] addr_remain3_3576;
address_decode_4 decoder_3_3576 = address_decode_4(addr_selector2_223[8],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3576,addr_remain3_3576);


wire[15:0] addr_selector3_3577;
wire[15:0] addr_remain3_3577;
address_decode_4 decoder_3_3577 = address_decode_4(addr_selector2_223[9],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3577,addr_remain3_3577);


wire[15:0] addr_selector3_3578;
wire[15:0] addr_remain3_3578;
address_decode_4 decoder_3_3578 = address_decode_4(addr_selector2_223[10],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3578,addr_remain3_3578);


wire[15:0] addr_selector3_3579;
wire[15:0] addr_remain3_3579;
address_decode_4 decoder_3_3579 = address_decode_4(addr_selector2_223[11],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3579,addr_remain3_3579);


wire[15:0] addr_selector3_3580;
wire[15:0] addr_remain3_3580;
address_decode_4 decoder_3_3580 = address_decode_4(addr_selector2_223[12],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3580,addr_remain3_3580);


wire[15:0] addr_selector3_3581;
wire[15:0] addr_remain3_3581;
address_decode_4 decoder_3_3581 = address_decode_4(addr_selector2_223[13],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3581,addr_remain3_3581);


wire[15:0] addr_selector3_3582;
wire[15:0] addr_remain3_3582;
address_decode_4 decoder_3_3582 = address_decode_4(addr_selector2_223[14],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3582,addr_remain3_3582);


wire[15:0] addr_selector3_3583;
wire[15:0] addr_remain3_3583;
address_decode_4 decoder_3_3583 = address_decode_4(addr_selector2_223[15],addr_remain2_223[15:0],addr_remain2_223,addr_selector3_3583,addr_remain3_3583);


wire[15:0] addr_selector3_3584;
wire[15:0] addr_remain3_3584;
address_decode_4 decoder_3_3584 = address_decode_4(addr_selector2_224[0],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3584,addr_remain3_3584);


wire[15:0] addr_selector3_3585;
wire[15:0] addr_remain3_3585;
address_decode_4 decoder_3_3585 = address_decode_4(addr_selector2_224[1],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3585,addr_remain3_3585);


wire[15:0] addr_selector3_3586;
wire[15:0] addr_remain3_3586;
address_decode_4 decoder_3_3586 = address_decode_4(addr_selector2_224[2],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3586,addr_remain3_3586);


wire[15:0] addr_selector3_3587;
wire[15:0] addr_remain3_3587;
address_decode_4 decoder_3_3587 = address_decode_4(addr_selector2_224[3],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3587,addr_remain3_3587);


wire[15:0] addr_selector3_3588;
wire[15:0] addr_remain3_3588;
address_decode_4 decoder_3_3588 = address_decode_4(addr_selector2_224[4],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3588,addr_remain3_3588);


wire[15:0] addr_selector3_3589;
wire[15:0] addr_remain3_3589;
address_decode_4 decoder_3_3589 = address_decode_4(addr_selector2_224[5],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3589,addr_remain3_3589);


wire[15:0] addr_selector3_3590;
wire[15:0] addr_remain3_3590;
address_decode_4 decoder_3_3590 = address_decode_4(addr_selector2_224[6],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3590,addr_remain3_3590);


wire[15:0] addr_selector3_3591;
wire[15:0] addr_remain3_3591;
address_decode_4 decoder_3_3591 = address_decode_4(addr_selector2_224[7],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3591,addr_remain3_3591);


wire[15:0] addr_selector3_3592;
wire[15:0] addr_remain3_3592;
address_decode_4 decoder_3_3592 = address_decode_4(addr_selector2_224[8],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3592,addr_remain3_3592);


wire[15:0] addr_selector3_3593;
wire[15:0] addr_remain3_3593;
address_decode_4 decoder_3_3593 = address_decode_4(addr_selector2_224[9],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3593,addr_remain3_3593);


wire[15:0] addr_selector3_3594;
wire[15:0] addr_remain3_3594;
address_decode_4 decoder_3_3594 = address_decode_4(addr_selector2_224[10],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3594,addr_remain3_3594);


wire[15:0] addr_selector3_3595;
wire[15:0] addr_remain3_3595;
address_decode_4 decoder_3_3595 = address_decode_4(addr_selector2_224[11],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3595,addr_remain3_3595);


wire[15:0] addr_selector3_3596;
wire[15:0] addr_remain3_3596;
address_decode_4 decoder_3_3596 = address_decode_4(addr_selector2_224[12],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3596,addr_remain3_3596);


wire[15:0] addr_selector3_3597;
wire[15:0] addr_remain3_3597;
address_decode_4 decoder_3_3597 = address_decode_4(addr_selector2_224[13],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3597,addr_remain3_3597);


wire[15:0] addr_selector3_3598;
wire[15:0] addr_remain3_3598;
address_decode_4 decoder_3_3598 = address_decode_4(addr_selector2_224[14],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3598,addr_remain3_3598);


wire[15:0] addr_selector3_3599;
wire[15:0] addr_remain3_3599;
address_decode_4 decoder_3_3599 = address_decode_4(addr_selector2_224[15],addr_remain2_224[15:0],addr_remain2_224,addr_selector3_3599,addr_remain3_3599);


wire[15:0] addr_selector3_3600;
wire[15:0] addr_remain3_3600;
address_decode_4 decoder_3_3600 = address_decode_4(addr_selector2_225[0],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3600,addr_remain3_3600);


wire[15:0] addr_selector3_3601;
wire[15:0] addr_remain3_3601;
address_decode_4 decoder_3_3601 = address_decode_4(addr_selector2_225[1],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3601,addr_remain3_3601);


wire[15:0] addr_selector3_3602;
wire[15:0] addr_remain3_3602;
address_decode_4 decoder_3_3602 = address_decode_4(addr_selector2_225[2],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3602,addr_remain3_3602);


wire[15:0] addr_selector3_3603;
wire[15:0] addr_remain3_3603;
address_decode_4 decoder_3_3603 = address_decode_4(addr_selector2_225[3],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3603,addr_remain3_3603);


wire[15:0] addr_selector3_3604;
wire[15:0] addr_remain3_3604;
address_decode_4 decoder_3_3604 = address_decode_4(addr_selector2_225[4],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3604,addr_remain3_3604);


wire[15:0] addr_selector3_3605;
wire[15:0] addr_remain3_3605;
address_decode_4 decoder_3_3605 = address_decode_4(addr_selector2_225[5],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3605,addr_remain3_3605);


wire[15:0] addr_selector3_3606;
wire[15:0] addr_remain3_3606;
address_decode_4 decoder_3_3606 = address_decode_4(addr_selector2_225[6],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3606,addr_remain3_3606);


wire[15:0] addr_selector3_3607;
wire[15:0] addr_remain3_3607;
address_decode_4 decoder_3_3607 = address_decode_4(addr_selector2_225[7],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3607,addr_remain3_3607);


wire[15:0] addr_selector3_3608;
wire[15:0] addr_remain3_3608;
address_decode_4 decoder_3_3608 = address_decode_4(addr_selector2_225[8],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3608,addr_remain3_3608);


wire[15:0] addr_selector3_3609;
wire[15:0] addr_remain3_3609;
address_decode_4 decoder_3_3609 = address_decode_4(addr_selector2_225[9],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3609,addr_remain3_3609);


wire[15:0] addr_selector3_3610;
wire[15:0] addr_remain3_3610;
address_decode_4 decoder_3_3610 = address_decode_4(addr_selector2_225[10],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3610,addr_remain3_3610);


wire[15:0] addr_selector3_3611;
wire[15:0] addr_remain3_3611;
address_decode_4 decoder_3_3611 = address_decode_4(addr_selector2_225[11],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3611,addr_remain3_3611);


wire[15:0] addr_selector3_3612;
wire[15:0] addr_remain3_3612;
address_decode_4 decoder_3_3612 = address_decode_4(addr_selector2_225[12],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3612,addr_remain3_3612);


wire[15:0] addr_selector3_3613;
wire[15:0] addr_remain3_3613;
address_decode_4 decoder_3_3613 = address_decode_4(addr_selector2_225[13],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3613,addr_remain3_3613);


wire[15:0] addr_selector3_3614;
wire[15:0] addr_remain3_3614;
address_decode_4 decoder_3_3614 = address_decode_4(addr_selector2_225[14],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3614,addr_remain3_3614);


wire[15:0] addr_selector3_3615;
wire[15:0] addr_remain3_3615;
address_decode_4 decoder_3_3615 = address_decode_4(addr_selector2_225[15],addr_remain2_225[15:0],addr_remain2_225,addr_selector3_3615,addr_remain3_3615);


wire[15:0] addr_selector3_3616;
wire[15:0] addr_remain3_3616;
address_decode_4 decoder_3_3616 = address_decode_4(addr_selector2_226[0],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3616,addr_remain3_3616);


wire[15:0] addr_selector3_3617;
wire[15:0] addr_remain3_3617;
address_decode_4 decoder_3_3617 = address_decode_4(addr_selector2_226[1],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3617,addr_remain3_3617);


wire[15:0] addr_selector3_3618;
wire[15:0] addr_remain3_3618;
address_decode_4 decoder_3_3618 = address_decode_4(addr_selector2_226[2],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3618,addr_remain3_3618);


wire[15:0] addr_selector3_3619;
wire[15:0] addr_remain3_3619;
address_decode_4 decoder_3_3619 = address_decode_4(addr_selector2_226[3],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3619,addr_remain3_3619);


wire[15:0] addr_selector3_3620;
wire[15:0] addr_remain3_3620;
address_decode_4 decoder_3_3620 = address_decode_4(addr_selector2_226[4],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3620,addr_remain3_3620);


wire[15:0] addr_selector3_3621;
wire[15:0] addr_remain3_3621;
address_decode_4 decoder_3_3621 = address_decode_4(addr_selector2_226[5],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3621,addr_remain3_3621);


wire[15:0] addr_selector3_3622;
wire[15:0] addr_remain3_3622;
address_decode_4 decoder_3_3622 = address_decode_4(addr_selector2_226[6],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3622,addr_remain3_3622);


wire[15:0] addr_selector3_3623;
wire[15:0] addr_remain3_3623;
address_decode_4 decoder_3_3623 = address_decode_4(addr_selector2_226[7],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3623,addr_remain3_3623);


wire[15:0] addr_selector3_3624;
wire[15:0] addr_remain3_3624;
address_decode_4 decoder_3_3624 = address_decode_4(addr_selector2_226[8],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3624,addr_remain3_3624);


wire[15:0] addr_selector3_3625;
wire[15:0] addr_remain3_3625;
address_decode_4 decoder_3_3625 = address_decode_4(addr_selector2_226[9],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3625,addr_remain3_3625);


wire[15:0] addr_selector3_3626;
wire[15:0] addr_remain3_3626;
address_decode_4 decoder_3_3626 = address_decode_4(addr_selector2_226[10],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3626,addr_remain3_3626);


wire[15:0] addr_selector3_3627;
wire[15:0] addr_remain3_3627;
address_decode_4 decoder_3_3627 = address_decode_4(addr_selector2_226[11],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3627,addr_remain3_3627);


wire[15:0] addr_selector3_3628;
wire[15:0] addr_remain3_3628;
address_decode_4 decoder_3_3628 = address_decode_4(addr_selector2_226[12],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3628,addr_remain3_3628);


wire[15:0] addr_selector3_3629;
wire[15:0] addr_remain3_3629;
address_decode_4 decoder_3_3629 = address_decode_4(addr_selector2_226[13],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3629,addr_remain3_3629);


wire[15:0] addr_selector3_3630;
wire[15:0] addr_remain3_3630;
address_decode_4 decoder_3_3630 = address_decode_4(addr_selector2_226[14],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3630,addr_remain3_3630);


wire[15:0] addr_selector3_3631;
wire[15:0] addr_remain3_3631;
address_decode_4 decoder_3_3631 = address_decode_4(addr_selector2_226[15],addr_remain2_226[15:0],addr_remain2_226,addr_selector3_3631,addr_remain3_3631);


wire[15:0] addr_selector3_3632;
wire[15:0] addr_remain3_3632;
address_decode_4 decoder_3_3632 = address_decode_4(addr_selector2_227[0],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3632,addr_remain3_3632);


wire[15:0] addr_selector3_3633;
wire[15:0] addr_remain3_3633;
address_decode_4 decoder_3_3633 = address_decode_4(addr_selector2_227[1],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3633,addr_remain3_3633);


wire[15:0] addr_selector3_3634;
wire[15:0] addr_remain3_3634;
address_decode_4 decoder_3_3634 = address_decode_4(addr_selector2_227[2],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3634,addr_remain3_3634);


wire[15:0] addr_selector3_3635;
wire[15:0] addr_remain3_3635;
address_decode_4 decoder_3_3635 = address_decode_4(addr_selector2_227[3],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3635,addr_remain3_3635);


wire[15:0] addr_selector3_3636;
wire[15:0] addr_remain3_3636;
address_decode_4 decoder_3_3636 = address_decode_4(addr_selector2_227[4],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3636,addr_remain3_3636);


wire[15:0] addr_selector3_3637;
wire[15:0] addr_remain3_3637;
address_decode_4 decoder_3_3637 = address_decode_4(addr_selector2_227[5],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3637,addr_remain3_3637);


wire[15:0] addr_selector3_3638;
wire[15:0] addr_remain3_3638;
address_decode_4 decoder_3_3638 = address_decode_4(addr_selector2_227[6],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3638,addr_remain3_3638);


wire[15:0] addr_selector3_3639;
wire[15:0] addr_remain3_3639;
address_decode_4 decoder_3_3639 = address_decode_4(addr_selector2_227[7],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3639,addr_remain3_3639);


wire[15:0] addr_selector3_3640;
wire[15:0] addr_remain3_3640;
address_decode_4 decoder_3_3640 = address_decode_4(addr_selector2_227[8],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3640,addr_remain3_3640);


wire[15:0] addr_selector3_3641;
wire[15:0] addr_remain3_3641;
address_decode_4 decoder_3_3641 = address_decode_4(addr_selector2_227[9],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3641,addr_remain3_3641);


wire[15:0] addr_selector3_3642;
wire[15:0] addr_remain3_3642;
address_decode_4 decoder_3_3642 = address_decode_4(addr_selector2_227[10],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3642,addr_remain3_3642);


wire[15:0] addr_selector3_3643;
wire[15:0] addr_remain3_3643;
address_decode_4 decoder_3_3643 = address_decode_4(addr_selector2_227[11],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3643,addr_remain3_3643);


wire[15:0] addr_selector3_3644;
wire[15:0] addr_remain3_3644;
address_decode_4 decoder_3_3644 = address_decode_4(addr_selector2_227[12],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3644,addr_remain3_3644);


wire[15:0] addr_selector3_3645;
wire[15:0] addr_remain3_3645;
address_decode_4 decoder_3_3645 = address_decode_4(addr_selector2_227[13],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3645,addr_remain3_3645);


wire[15:0] addr_selector3_3646;
wire[15:0] addr_remain3_3646;
address_decode_4 decoder_3_3646 = address_decode_4(addr_selector2_227[14],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3646,addr_remain3_3646);


wire[15:0] addr_selector3_3647;
wire[15:0] addr_remain3_3647;
address_decode_4 decoder_3_3647 = address_decode_4(addr_selector2_227[15],addr_remain2_227[15:0],addr_remain2_227,addr_selector3_3647,addr_remain3_3647);


wire[15:0] addr_selector3_3648;
wire[15:0] addr_remain3_3648;
address_decode_4 decoder_3_3648 = address_decode_4(addr_selector2_228[0],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3648,addr_remain3_3648);


wire[15:0] addr_selector3_3649;
wire[15:0] addr_remain3_3649;
address_decode_4 decoder_3_3649 = address_decode_4(addr_selector2_228[1],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3649,addr_remain3_3649);


wire[15:0] addr_selector3_3650;
wire[15:0] addr_remain3_3650;
address_decode_4 decoder_3_3650 = address_decode_4(addr_selector2_228[2],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3650,addr_remain3_3650);


wire[15:0] addr_selector3_3651;
wire[15:0] addr_remain3_3651;
address_decode_4 decoder_3_3651 = address_decode_4(addr_selector2_228[3],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3651,addr_remain3_3651);


wire[15:0] addr_selector3_3652;
wire[15:0] addr_remain3_3652;
address_decode_4 decoder_3_3652 = address_decode_4(addr_selector2_228[4],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3652,addr_remain3_3652);


wire[15:0] addr_selector3_3653;
wire[15:0] addr_remain3_3653;
address_decode_4 decoder_3_3653 = address_decode_4(addr_selector2_228[5],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3653,addr_remain3_3653);


wire[15:0] addr_selector3_3654;
wire[15:0] addr_remain3_3654;
address_decode_4 decoder_3_3654 = address_decode_4(addr_selector2_228[6],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3654,addr_remain3_3654);


wire[15:0] addr_selector3_3655;
wire[15:0] addr_remain3_3655;
address_decode_4 decoder_3_3655 = address_decode_4(addr_selector2_228[7],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3655,addr_remain3_3655);


wire[15:0] addr_selector3_3656;
wire[15:0] addr_remain3_3656;
address_decode_4 decoder_3_3656 = address_decode_4(addr_selector2_228[8],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3656,addr_remain3_3656);


wire[15:0] addr_selector3_3657;
wire[15:0] addr_remain3_3657;
address_decode_4 decoder_3_3657 = address_decode_4(addr_selector2_228[9],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3657,addr_remain3_3657);


wire[15:0] addr_selector3_3658;
wire[15:0] addr_remain3_3658;
address_decode_4 decoder_3_3658 = address_decode_4(addr_selector2_228[10],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3658,addr_remain3_3658);


wire[15:0] addr_selector3_3659;
wire[15:0] addr_remain3_3659;
address_decode_4 decoder_3_3659 = address_decode_4(addr_selector2_228[11],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3659,addr_remain3_3659);


wire[15:0] addr_selector3_3660;
wire[15:0] addr_remain3_3660;
address_decode_4 decoder_3_3660 = address_decode_4(addr_selector2_228[12],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3660,addr_remain3_3660);


wire[15:0] addr_selector3_3661;
wire[15:0] addr_remain3_3661;
address_decode_4 decoder_3_3661 = address_decode_4(addr_selector2_228[13],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3661,addr_remain3_3661);


wire[15:0] addr_selector3_3662;
wire[15:0] addr_remain3_3662;
address_decode_4 decoder_3_3662 = address_decode_4(addr_selector2_228[14],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3662,addr_remain3_3662);


wire[15:0] addr_selector3_3663;
wire[15:0] addr_remain3_3663;
address_decode_4 decoder_3_3663 = address_decode_4(addr_selector2_228[15],addr_remain2_228[15:0],addr_remain2_228,addr_selector3_3663,addr_remain3_3663);


wire[15:0] addr_selector3_3664;
wire[15:0] addr_remain3_3664;
address_decode_4 decoder_3_3664 = address_decode_4(addr_selector2_229[0],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3664,addr_remain3_3664);


wire[15:0] addr_selector3_3665;
wire[15:0] addr_remain3_3665;
address_decode_4 decoder_3_3665 = address_decode_4(addr_selector2_229[1],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3665,addr_remain3_3665);


wire[15:0] addr_selector3_3666;
wire[15:0] addr_remain3_3666;
address_decode_4 decoder_3_3666 = address_decode_4(addr_selector2_229[2],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3666,addr_remain3_3666);


wire[15:0] addr_selector3_3667;
wire[15:0] addr_remain3_3667;
address_decode_4 decoder_3_3667 = address_decode_4(addr_selector2_229[3],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3667,addr_remain3_3667);


wire[15:0] addr_selector3_3668;
wire[15:0] addr_remain3_3668;
address_decode_4 decoder_3_3668 = address_decode_4(addr_selector2_229[4],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3668,addr_remain3_3668);


wire[15:0] addr_selector3_3669;
wire[15:0] addr_remain3_3669;
address_decode_4 decoder_3_3669 = address_decode_4(addr_selector2_229[5],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3669,addr_remain3_3669);


wire[15:0] addr_selector3_3670;
wire[15:0] addr_remain3_3670;
address_decode_4 decoder_3_3670 = address_decode_4(addr_selector2_229[6],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3670,addr_remain3_3670);


wire[15:0] addr_selector3_3671;
wire[15:0] addr_remain3_3671;
address_decode_4 decoder_3_3671 = address_decode_4(addr_selector2_229[7],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3671,addr_remain3_3671);


wire[15:0] addr_selector3_3672;
wire[15:0] addr_remain3_3672;
address_decode_4 decoder_3_3672 = address_decode_4(addr_selector2_229[8],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3672,addr_remain3_3672);


wire[15:0] addr_selector3_3673;
wire[15:0] addr_remain3_3673;
address_decode_4 decoder_3_3673 = address_decode_4(addr_selector2_229[9],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3673,addr_remain3_3673);


wire[15:0] addr_selector3_3674;
wire[15:0] addr_remain3_3674;
address_decode_4 decoder_3_3674 = address_decode_4(addr_selector2_229[10],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3674,addr_remain3_3674);


wire[15:0] addr_selector3_3675;
wire[15:0] addr_remain3_3675;
address_decode_4 decoder_3_3675 = address_decode_4(addr_selector2_229[11],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3675,addr_remain3_3675);


wire[15:0] addr_selector3_3676;
wire[15:0] addr_remain3_3676;
address_decode_4 decoder_3_3676 = address_decode_4(addr_selector2_229[12],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3676,addr_remain3_3676);


wire[15:0] addr_selector3_3677;
wire[15:0] addr_remain3_3677;
address_decode_4 decoder_3_3677 = address_decode_4(addr_selector2_229[13],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3677,addr_remain3_3677);


wire[15:0] addr_selector3_3678;
wire[15:0] addr_remain3_3678;
address_decode_4 decoder_3_3678 = address_decode_4(addr_selector2_229[14],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3678,addr_remain3_3678);


wire[15:0] addr_selector3_3679;
wire[15:0] addr_remain3_3679;
address_decode_4 decoder_3_3679 = address_decode_4(addr_selector2_229[15],addr_remain2_229[15:0],addr_remain2_229,addr_selector3_3679,addr_remain3_3679);


wire[15:0] addr_selector3_3680;
wire[15:0] addr_remain3_3680;
address_decode_4 decoder_3_3680 = address_decode_4(addr_selector2_230[0],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3680,addr_remain3_3680);


wire[15:0] addr_selector3_3681;
wire[15:0] addr_remain3_3681;
address_decode_4 decoder_3_3681 = address_decode_4(addr_selector2_230[1],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3681,addr_remain3_3681);


wire[15:0] addr_selector3_3682;
wire[15:0] addr_remain3_3682;
address_decode_4 decoder_3_3682 = address_decode_4(addr_selector2_230[2],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3682,addr_remain3_3682);


wire[15:0] addr_selector3_3683;
wire[15:0] addr_remain3_3683;
address_decode_4 decoder_3_3683 = address_decode_4(addr_selector2_230[3],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3683,addr_remain3_3683);


wire[15:0] addr_selector3_3684;
wire[15:0] addr_remain3_3684;
address_decode_4 decoder_3_3684 = address_decode_4(addr_selector2_230[4],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3684,addr_remain3_3684);


wire[15:0] addr_selector3_3685;
wire[15:0] addr_remain3_3685;
address_decode_4 decoder_3_3685 = address_decode_4(addr_selector2_230[5],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3685,addr_remain3_3685);


wire[15:0] addr_selector3_3686;
wire[15:0] addr_remain3_3686;
address_decode_4 decoder_3_3686 = address_decode_4(addr_selector2_230[6],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3686,addr_remain3_3686);


wire[15:0] addr_selector3_3687;
wire[15:0] addr_remain3_3687;
address_decode_4 decoder_3_3687 = address_decode_4(addr_selector2_230[7],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3687,addr_remain3_3687);


wire[15:0] addr_selector3_3688;
wire[15:0] addr_remain3_3688;
address_decode_4 decoder_3_3688 = address_decode_4(addr_selector2_230[8],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3688,addr_remain3_3688);


wire[15:0] addr_selector3_3689;
wire[15:0] addr_remain3_3689;
address_decode_4 decoder_3_3689 = address_decode_4(addr_selector2_230[9],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3689,addr_remain3_3689);


wire[15:0] addr_selector3_3690;
wire[15:0] addr_remain3_3690;
address_decode_4 decoder_3_3690 = address_decode_4(addr_selector2_230[10],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3690,addr_remain3_3690);


wire[15:0] addr_selector3_3691;
wire[15:0] addr_remain3_3691;
address_decode_4 decoder_3_3691 = address_decode_4(addr_selector2_230[11],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3691,addr_remain3_3691);


wire[15:0] addr_selector3_3692;
wire[15:0] addr_remain3_3692;
address_decode_4 decoder_3_3692 = address_decode_4(addr_selector2_230[12],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3692,addr_remain3_3692);


wire[15:0] addr_selector3_3693;
wire[15:0] addr_remain3_3693;
address_decode_4 decoder_3_3693 = address_decode_4(addr_selector2_230[13],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3693,addr_remain3_3693);


wire[15:0] addr_selector3_3694;
wire[15:0] addr_remain3_3694;
address_decode_4 decoder_3_3694 = address_decode_4(addr_selector2_230[14],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3694,addr_remain3_3694);


wire[15:0] addr_selector3_3695;
wire[15:0] addr_remain3_3695;
address_decode_4 decoder_3_3695 = address_decode_4(addr_selector2_230[15],addr_remain2_230[15:0],addr_remain2_230,addr_selector3_3695,addr_remain3_3695);


wire[15:0] addr_selector3_3696;
wire[15:0] addr_remain3_3696;
address_decode_4 decoder_3_3696 = address_decode_4(addr_selector2_231[0],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3696,addr_remain3_3696);


wire[15:0] addr_selector3_3697;
wire[15:0] addr_remain3_3697;
address_decode_4 decoder_3_3697 = address_decode_4(addr_selector2_231[1],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3697,addr_remain3_3697);


wire[15:0] addr_selector3_3698;
wire[15:0] addr_remain3_3698;
address_decode_4 decoder_3_3698 = address_decode_4(addr_selector2_231[2],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3698,addr_remain3_3698);


wire[15:0] addr_selector3_3699;
wire[15:0] addr_remain3_3699;
address_decode_4 decoder_3_3699 = address_decode_4(addr_selector2_231[3],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3699,addr_remain3_3699);


wire[15:0] addr_selector3_3700;
wire[15:0] addr_remain3_3700;
address_decode_4 decoder_3_3700 = address_decode_4(addr_selector2_231[4],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3700,addr_remain3_3700);


wire[15:0] addr_selector3_3701;
wire[15:0] addr_remain3_3701;
address_decode_4 decoder_3_3701 = address_decode_4(addr_selector2_231[5],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3701,addr_remain3_3701);


wire[15:0] addr_selector3_3702;
wire[15:0] addr_remain3_3702;
address_decode_4 decoder_3_3702 = address_decode_4(addr_selector2_231[6],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3702,addr_remain3_3702);


wire[15:0] addr_selector3_3703;
wire[15:0] addr_remain3_3703;
address_decode_4 decoder_3_3703 = address_decode_4(addr_selector2_231[7],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3703,addr_remain3_3703);


wire[15:0] addr_selector3_3704;
wire[15:0] addr_remain3_3704;
address_decode_4 decoder_3_3704 = address_decode_4(addr_selector2_231[8],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3704,addr_remain3_3704);


wire[15:0] addr_selector3_3705;
wire[15:0] addr_remain3_3705;
address_decode_4 decoder_3_3705 = address_decode_4(addr_selector2_231[9],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3705,addr_remain3_3705);


wire[15:0] addr_selector3_3706;
wire[15:0] addr_remain3_3706;
address_decode_4 decoder_3_3706 = address_decode_4(addr_selector2_231[10],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3706,addr_remain3_3706);


wire[15:0] addr_selector3_3707;
wire[15:0] addr_remain3_3707;
address_decode_4 decoder_3_3707 = address_decode_4(addr_selector2_231[11],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3707,addr_remain3_3707);


wire[15:0] addr_selector3_3708;
wire[15:0] addr_remain3_3708;
address_decode_4 decoder_3_3708 = address_decode_4(addr_selector2_231[12],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3708,addr_remain3_3708);


wire[15:0] addr_selector3_3709;
wire[15:0] addr_remain3_3709;
address_decode_4 decoder_3_3709 = address_decode_4(addr_selector2_231[13],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3709,addr_remain3_3709);


wire[15:0] addr_selector3_3710;
wire[15:0] addr_remain3_3710;
address_decode_4 decoder_3_3710 = address_decode_4(addr_selector2_231[14],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3710,addr_remain3_3710);


wire[15:0] addr_selector3_3711;
wire[15:0] addr_remain3_3711;
address_decode_4 decoder_3_3711 = address_decode_4(addr_selector2_231[15],addr_remain2_231[15:0],addr_remain2_231,addr_selector3_3711,addr_remain3_3711);


wire[15:0] addr_selector3_3712;
wire[15:0] addr_remain3_3712;
address_decode_4 decoder_3_3712 = address_decode_4(addr_selector2_232[0],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3712,addr_remain3_3712);


wire[15:0] addr_selector3_3713;
wire[15:0] addr_remain3_3713;
address_decode_4 decoder_3_3713 = address_decode_4(addr_selector2_232[1],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3713,addr_remain3_3713);


wire[15:0] addr_selector3_3714;
wire[15:0] addr_remain3_3714;
address_decode_4 decoder_3_3714 = address_decode_4(addr_selector2_232[2],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3714,addr_remain3_3714);


wire[15:0] addr_selector3_3715;
wire[15:0] addr_remain3_3715;
address_decode_4 decoder_3_3715 = address_decode_4(addr_selector2_232[3],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3715,addr_remain3_3715);


wire[15:0] addr_selector3_3716;
wire[15:0] addr_remain3_3716;
address_decode_4 decoder_3_3716 = address_decode_4(addr_selector2_232[4],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3716,addr_remain3_3716);


wire[15:0] addr_selector3_3717;
wire[15:0] addr_remain3_3717;
address_decode_4 decoder_3_3717 = address_decode_4(addr_selector2_232[5],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3717,addr_remain3_3717);


wire[15:0] addr_selector3_3718;
wire[15:0] addr_remain3_3718;
address_decode_4 decoder_3_3718 = address_decode_4(addr_selector2_232[6],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3718,addr_remain3_3718);


wire[15:0] addr_selector3_3719;
wire[15:0] addr_remain3_3719;
address_decode_4 decoder_3_3719 = address_decode_4(addr_selector2_232[7],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3719,addr_remain3_3719);


wire[15:0] addr_selector3_3720;
wire[15:0] addr_remain3_3720;
address_decode_4 decoder_3_3720 = address_decode_4(addr_selector2_232[8],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3720,addr_remain3_3720);


wire[15:0] addr_selector3_3721;
wire[15:0] addr_remain3_3721;
address_decode_4 decoder_3_3721 = address_decode_4(addr_selector2_232[9],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3721,addr_remain3_3721);


wire[15:0] addr_selector3_3722;
wire[15:0] addr_remain3_3722;
address_decode_4 decoder_3_3722 = address_decode_4(addr_selector2_232[10],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3722,addr_remain3_3722);


wire[15:0] addr_selector3_3723;
wire[15:0] addr_remain3_3723;
address_decode_4 decoder_3_3723 = address_decode_4(addr_selector2_232[11],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3723,addr_remain3_3723);


wire[15:0] addr_selector3_3724;
wire[15:0] addr_remain3_3724;
address_decode_4 decoder_3_3724 = address_decode_4(addr_selector2_232[12],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3724,addr_remain3_3724);


wire[15:0] addr_selector3_3725;
wire[15:0] addr_remain3_3725;
address_decode_4 decoder_3_3725 = address_decode_4(addr_selector2_232[13],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3725,addr_remain3_3725);


wire[15:0] addr_selector3_3726;
wire[15:0] addr_remain3_3726;
address_decode_4 decoder_3_3726 = address_decode_4(addr_selector2_232[14],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3726,addr_remain3_3726);


wire[15:0] addr_selector3_3727;
wire[15:0] addr_remain3_3727;
address_decode_4 decoder_3_3727 = address_decode_4(addr_selector2_232[15],addr_remain2_232[15:0],addr_remain2_232,addr_selector3_3727,addr_remain3_3727);


wire[15:0] addr_selector3_3728;
wire[15:0] addr_remain3_3728;
address_decode_4 decoder_3_3728 = address_decode_4(addr_selector2_233[0],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3728,addr_remain3_3728);


wire[15:0] addr_selector3_3729;
wire[15:0] addr_remain3_3729;
address_decode_4 decoder_3_3729 = address_decode_4(addr_selector2_233[1],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3729,addr_remain3_3729);


wire[15:0] addr_selector3_3730;
wire[15:0] addr_remain3_3730;
address_decode_4 decoder_3_3730 = address_decode_4(addr_selector2_233[2],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3730,addr_remain3_3730);


wire[15:0] addr_selector3_3731;
wire[15:0] addr_remain3_3731;
address_decode_4 decoder_3_3731 = address_decode_4(addr_selector2_233[3],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3731,addr_remain3_3731);


wire[15:0] addr_selector3_3732;
wire[15:0] addr_remain3_3732;
address_decode_4 decoder_3_3732 = address_decode_4(addr_selector2_233[4],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3732,addr_remain3_3732);


wire[15:0] addr_selector3_3733;
wire[15:0] addr_remain3_3733;
address_decode_4 decoder_3_3733 = address_decode_4(addr_selector2_233[5],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3733,addr_remain3_3733);


wire[15:0] addr_selector3_3734;
wire[15:0] addr_remain3_3734;
address_decode_4 decoder_3_3734 = address_decode_4(addr_selector2_233[6],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3734,addr_remain3_3734);


wire[15:0] addr_selector3_3735;
wire[15:0] addr_remain3_3735;
address_decode_4 decoder_3_3735 = address_decode_4(addr_selector2_233[7],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3735,addr_remain3_3735);


wire[15:0] addr_selector3_3736;
wire[15:0] addr_remain3_3736;
address_decode_4 decoder_3_3736 = address_decode_4(addr_selector2_233[8],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3736,addr_remain3_3736);


wire[15:0] addr_selector3_3737;
wire[15:0] addr_remain3_3737;
address_decode_4 decoder_3_3737 = address_decode_4(addr_selector2_233[9],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3737,addr_remain3_3737);


wire[15:0] addr_selector3_3738;
wire[15:0] addr_remain3_3738;
address_decode_4 decoder_3_3738 = address_decode_4(addr_selector2_233[10],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3738,addr_remain3_3738);


wire[15:0] addr_selector3_3739;
wire[15:0] addr_remain3_3739;
address_decode_4 decoder_3_3739 = address_decode_4(addr_selector2_233[11],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3739,addr_remain3_3739);


wire[15:0] addr_selector3_3740;
wire[15:0] addr_remain3_3740;
address_decode_4 decoder_3_3740 = address_decode_4(addr_selector2_233[12],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3740,addr_remain3_3740);


wire[15:0] addr_selector3_3741;
wire[15:0] addr_remain3_3741;
address_decode_4 decoder_3_3741 = address_decode_4(addr_selector2_233[13],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3741,addr_remain3_3741);


wire[15:0] addr_selector3_3742;
wire[15:0] addr_remain3_3742;
address_decode_4 decoder_3_3742 = address_decode_4(addr_selector2_233[14],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3742,addr_remain3_3742);


wire[15:0] addr_selector3_3743;
wire[15:0] addr_remain3_3743;
address_decode_4 decoder_3_3743 = address_decode_4(addr_selector2_233[15],addr_remain2_233[15:0],addr_remain2_233,addr_selector3_3743,addr_remain3_3743);


wire[15:0] addr_selector3_3744;
wire[15:0] addr_remain3_3744;
address_decode_4 decoder_3_3744 = address_decode_4(addr_selector2_234[0],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3744,addr_remain3_3744);


wire[15:0] addr_selector3_3745;
wire[15:0] addr_remain3_3745;
address_decode_4 decoder_3_3745 = address_decode_4(addr_selector2_234[1],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3745,addr_remain3_3745);


wire[15:0] addr_selector3_3746;
wire[15:0] addr_remain3_3746;
address_decode_4 decoder_3_3746 = address_decode_4(addr_selector2_234[2],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3746,addr_remain3_3746);


wire[15:0] addr_selector3_3747;
wire[15:0] addr_remain3_3747;
address_decode_4 decoder_3_3747 = address_decode_4(addr_selector2_234[3],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3747,addr_remain3_3747);


wire[15:0] addr_selector3_3748;
wire[15:0] addr_remain3_3748;
address_decode_4 decoder_3_3748 = address_decode_4(addr_selector2_234[4],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3748,addr_remain3_3748);


wire[15:0] addr_selector3_3749;
wire[15:0] addr_remain3_3749;
address_decode_4 decoder_3_3749 = address_decode_4(addr_selector2_234[5],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3749,addr_remain3_3749);


wire[15:0] addr_selector3_3750;
wire[15:0] addr_remain3_3750;
address_decode_4 decoder_3_3750 = address_decode_4(addr_selector2_234[6],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3750,addr_remain3_3750);


wire[15:0] addr_selector3_3751;
wire[15:0] addr_remain3_3751;
address_decode_4 decoder_3_3751 = address_decode_4(addr_selector2_234[7],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3751,addr_remain3_3751);


wire[15:0] addr_selector3_3752;
wire[15:0] addr_remain3_3752;
address_decode_4 decoder_3_3752 = address_decode_4(addr_selector2_234[8],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3752,addr_remain3_3752);


wire[15:0] addr_selector3_3753;
wire[15:0] addr_remain3_3753;
address_decode_4 decoder_3_3753 = address_decode_4(addr_selector2_234[9],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3753,addr_remain3_3753);


wire[15:0] addr_selector3_3754;
wire[15:0] addr_remain3_3754;
address_decode_4 decoder_3_3754 = address_decode_4(addr_selector2_234[10],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3754,addr_remain3_3754);


wire[15:0] addr_selector3_3755;
wire[15:0] addr_remain3_3755;
address_decode_4 decoder_3_3755 = address_decode_4(addr_selector2_234[11],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3755,addr_remain3_3755);


wire[15:0] addr_selector3_3756;
wire[15:0] addr_remain3_3756;
address_decode_4 decoder_3_3756 = address_decode_4(addr_selector2_234[12],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3756,addr_remain3_3756);


wire[15:0] addr_selector3_3757;
wire[15:0] addr_remain3_3757;
address_decode_4 decoder_3_3757 = address_decode_4(addr_selector2_234[13],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3757,addr_remain3_3757);


wire[15:0] addr_selector3_3758;
wire[15:0] addr_remain3_3758;
address_decode_4 decoder_3_3758 = address_decode_4(addr_selector2_234[14],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3758,addr_remain3_3758);


wire[15:0] addr_selector3_3759;
wire[15:0] addr_remain3_3759;
address_decode_4 decoder_3_3759 = address_decode_4(addr_selector2_234[15],addr_remain2_234[15:0],addr_remain2_234,addr_selector3_3759,addr_remain3_3759);


wire[15:0] addr_selector3_3760;
wire[15:0] addr_remain3_3760;
address_decode_4 decoder_3_3760 = address_decode_4(addr_selector2_235[0],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3760,addr_remain3_3760);


wire[15:0] addr_selector3_3761;
wire[15:0] addr_remain3_3761;
address_decode_4 decoder_3_3761 = address_decode_4(addr_selector2_235[1],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3761,addr_remain3_3761);


wire[15:0] addr_selector3_3762;
wire[15:0] addr_remain3_3762;
address_decode_4 decoder_3_3762 = address_decode_4(addr_selector2_235[2],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3762,addr_remain3_3762);


wire[15:0] addr_selector3_3763;
wire[15:0] addr_remain3_3763;
address_decode_4 decoder_3_3763 = address_decode_4(addr_selector2_235[3],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3763,addr_remain3_3763);


wire[15:0] addr_selector3_3764;
wire[15:0] addr_remain3_3764;
address_decode_4 decoder_3_3764 = address_decode_4(addr_selector2_235[4],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3764,addr_remain3_3764);


wire[15:0] addr_selector3_3765;
wire[15:0] addr_remain3_3765;
address_decode_4 decoder_3_3765 = address_decode_4(addr_selector2_235[5],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3765,addr_remain3_3765);


wire[15:0] addr_selector3_3766;
wire[15:0] addr_remain3_3766;
address_decode_4 decoder_3_3766 = address_decode_4(addr_selector2_235[6],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3766,addr_remain3_3766);


wire[15:0] addr_selector3_3767;
wire[15:0] addr_remain3_3767;
address_decode_4 decoder_3_3767 = address_decode_4(addr_selector2_235[7],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3767,addr_remain3_3767);


wire[15:0] addr_selector3_3768;
wire[15:0] addr_remain3_3768;
address_decode_4 decoder_3_3768 = address_decode_4(addr_selector2_235[8],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3768,addr_remain3_3768);


wire[15:0] addr_selector3_3769;
wire[15:0] addr_remain3_3769;
address_decode_4 decoder_3_3769 = address_decode_4(addr_selector2_235[9],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3769,addr_remain3_3769);


wire[15:0] addr_selector3_3770;
wire[15:0] addr_remain3_3770;
address_decode_4 decoder_3_3770 = address_decode_4(addr_selector2_235[10],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3770,addr_remain3_3770);


wire[15:0] addr_selector3_3771;
wire[15:0] addr_remain3_3771;
address_decode_4 decoder_3_3771 = address_decode_4(addr_selector2_235[11],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3771,addr_remain3_3771);


wire[15:0] addr_selector3_3772;
wire[15:0] addr_remain3_3772;
address_decode_4 decoder_3_3772 = address_decode_4(addr_selector2_235[12],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3772,addr_remain3_3772);


wire[15:0] addr_selector3_3773;
wire[15:0] addr_remain3_3773;
address_decode_4 decoder_3_3773 = address_decode_4(addr_selector2_235[13],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3773,addr_remain3_3773);


wire[15:0] addr_selector3_3774;
wire[15:0] addr_remain3_3774;
address_decode_4 decoder_3_3774 = address_decode_4(addr_selector2_235[14],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3774,addr_remain3_3774);


wire[15:0] addr_selector3_3775;
wire[15:0] addr_remain3_3775;
address_decode_4 decoder_3_3775 = address_decode_4(addr_selector2_235[15],addr_remain2_235[15:0],addr_remain2_235,addr_selector3_3775,addr_remain3_3775);


wire[15:0] addr_selector3_3776;
wire[15:0] addr_remain3_3776;
address_decode_4 decoder_3_3776 = address_decode_4(addr_selector2_236[0],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3776,addr_remain3_3776);


wire[15:0] addr_selector3_3777;
wire[15:0] addr_remain3_3777;
address_decode_4 decoder_3_3777 = address_decode_4(addr_selector2_236[1],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3777,addr_remain3_3777);


wire[15:0] addr_selector3_3778;
wire[15:0] addr_remain3_3778;
address_decode_4 decoder_3_3778 = address_decode_4(addr_selector2_236[2],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3778,addr_remain3_3778);


wire[15:0] addr_selector3_3779;
wire[15:0] addr_remain3_3779;
address_decode_4 decoder_3_3779 = address_decode_4(addr_selector2_236[3],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3779,addr_remain3_3779);


wire[15:0] addr_selector3_3780;
wire[15:0] addr_remain3_3780;
address_decode_4 decoder_3_3780 = address_decode_4(addr_selector2_236[4],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3780,addr_remain3_3780);


wire[15:0] addr_selector3_3781;
wire[15:0] addr_remain3_3781;
address_decode_4 decoder_3_3781 = address_decode_4(addr_selector2_236[5],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3781,addr_remain3_3781);


wire[15:0] addr_selector3_3782;
wire[15:0] addr_remain3_3782;
address_decode_4 decoder_3_3782 = address_decode_4(addr_selector2_236[6],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3782,addr_remain3_3782);


wire[15:0] addr_selector3_3783;
wire[15:0] addr_remain3_3783;
address_decode_4 decoder_3_3783 = address_decode_4(addr_selector2_236[7],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3783,addr_remain3_3783);


wire[15:0] addr_selector3_3784;
wire[15:0] addr_remain3_3784;
address_decode_4 decoder_3_3784 = address_decode_4(addr_selector2_236[8],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3784,addr_remain3_3784);


wire[15:0] addr_selector3_3785;
wire[15:0] addr_remain3_3785;
address_decode_4 decoder_3_3785 = address_decode_4(addr_selector2_236[9],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3785,addr_remain3_3785);


wire[15:0] addr_selector3_3786;
wire[15:0] addr_remain3_3786;
address_decode_4 decoder_3_3786 = address_decode_4(addr_selector2_236[10],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3786,addr_remain3_3786);


wire[15:0] addr_selector3_3787;
wire[15:0] addr_remain3_3787;
address_decode_4 decoder_3_3787 = address_decode_4(addr_selector2_236[11],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3787,addr_remain3_3787);


wire[15:0] addr_selector3_3788;
wire[15:0] addr_remain3_3788;
address_decode_4 decoder_3_3788 = address_decode_4(addr_selector2_236[12],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3788,addr_remain3_3788);


wire[15:0] addr_selector3_3789;
wire[15:0] addr_remain3_3789;
address_decode_4 decoder_3_3789 = address_decode_4(addr_selector2_236[13],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3789,addr_remain3_3789);


wire[15:0] addr_selector3_3790;
wire[15:0] addr_remain3_3790;
address_decode_4 decoder_3_3790 = address_decode_4(addr_selector2_236[14],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3790,addr_remain3_3790);


wire[15:0] addr_selector3_3791;
wire[15:0] addr_remain3_3791;
address_decode_4 decoder_3_3791 = address_decode_4(addr_selector2_236[15],addr_remain2_236[15:0],addr_remain2_236,addr_selector3_3791,addr_remain3_3791);


wire[15:0] addr_selector3_3792;
wire[15:0] addr_remain3_3792;
address_decode_4 decoder_3_3792 = address_decode_4(addr_selector2_237[0],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3792,addr_remain3_3792);


wire[15:0] addr_selector3_3793;
wire[15:0] addr_remain3_3793;
address_decode_4 decoder_3_3793 = address_decode_4(addr_selector2_237[1],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3793,addr_remain3_3793);


wire[15:0] addr_selector3_3794;
wire[15:0] addr_remain3_3794;
address_decode_4 decoder_3_3794 = address_decode_4(addr_selector2_237[2],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3794,addr_remain3_3794);


wire[15:0] addr_selector3_3795;
wire[15:0] addr_remain3_3795;
address_decode_4 decoder_3_3795 = address_decode_4(addr_selector2_237[3],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3795,addr_remain3_3795);


wire[15:0] addr_selector3_3796;
wire[15:0] addr_remain3_3796;
address_decode_4 decoder_3_3796 = address_decode_4(addr_selector2_237[4],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3796,addr_remain3_3796);


wire[15:0] addr_selector3_3797;
wire[15:0] addr_remain3_3797;
address_decode_4 decoder_3_3797 = address_decode_4(addr_selector2_237[5],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3797,addr_remain3_3797);


wire[15:0] addr_selector3_3798;
wire[15:0] addr_remain3_3798;
address_decode_4 decoder_3_3798 = address_decode_4(addr_selector2_237[6],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3798,addr_remain3_3798);


wire[15:0] addr_selector3_3799;
wire[15:0] addr_remain3_3799;
address_decode_4 decoder_3_3799 = address_decode_4(addr_selector2_237[7],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3799,addr_remain3_3799);


wire[15:0] addr_selector3_3800;
wire[15:0] addr_remain3_3800;
address_decode_4 decoder_3_3800 = address_decode_4(addr_selector2_237[8],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3800,addr_remain3_3800);


wire[15:0] addr_selector3_3801;
wire[15:0] addr_remain3_3801;
address_decode_4 decoder_3_3801 = address_decode_4(addr_selector2_237[9],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3801,addr_remain3_3801);


wire[15:0] addr_selector3_3802;
wire[15:0] addr_remain3_3802;
address_decode_4 decoder_3_3802 = address_decode_4(addr_selector2_237[10],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3802,addr_remain3_3802);


wire[15:0] addr_selector3_3803;
wire[15:0] addr_remain3_3803;
address_decode_4 decoder_3_3803 = address_decode_4(addr_selector2_237[11],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3803,addr_remain3_3803);


wire[15:0] addr_selector3_3804;
wire[15:0] addr_remain3_3804;
address_decode_4 decoder_3_3804 = address_decode_4(addr_selector2_237[12],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3804,addr_remain3_3804);


wire[15:0] addr_selector3_3805;
wire[15:0] addr_remain3_3805;
address_decode_4 decoder_3_3805 = address_decode_4(addr_selector2_237[13],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3805,addr_remain3_3805);


wire[15:0] addr_selector3_3806;
wire[15:0] addr_remain3_3806;
address_decode_4 decoder_3_3806 = address_decode_4(addr_selector2_237[14],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3806,addr_remain3_3806);


wire[15:0] addr_selector3_3807;
wire[15:0] addr_remain3_3807;
address_decode_4 decoder_3_3807 = address_decode_4(addr_selector2_237[15],addr_remain2_237[15:0],addr_remain2_237,addr_selector3_3807,addr_remain3_3807);


wire[15:0] addr_selector3_3808;
wire[15:0] addr_remain3_3808;
address_decode_4 decoder_3_3808 = address_decode_4(addr_selector2_238[0],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3808,addr_remain3_3808);


wire[15:0] addr_selector3_3809;
wire[15:0] addr_remain3_3809;
address_decode_4 decoder_3_3809 = address_decode_4(addr_selector2_238[1],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3809,addr_remain3_3809);


wire[15:0] addr_selector3_3810;
wire[15:0] addr_remain3_3810;
address_decode_4 decoder_3_3810 = address_decode_4(addr_selector2_238[2],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3810,addr_remain3_3810);


wire[15:0] addr_selector3_3811;
wire[15:0] addr_remain3_3811;
address_decode_4 decoder_3_3811 = address_decode_4(addr_selector2_238[3],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3811,addr_remain3_3811);


wire[15:0] addr_selector3_3812;
wire[15:0] addr_remain3_3812;
address_decode_4 decoder_3_3812 = address_decode_4(addr_selector2_238[4],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3812,addr_remain3_3812);


wire[15:0] addr_selector3_3813;
wire[15:0] addr_remain3_3813;
address_decode_4 decoder_3_3813 = address_decode_4(addr_selector2_238[5],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3813,addr_remain3_3813);


wire[15:0] addr_selector3_3814;
wire[15:0] addr_remain3_3814;
address_decode_4 decoder_3_3814 = address_decode_4(addr_selector2_238[6],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3814,addr_remain3_3814);


wire[15:0] addr_selector3_3815;
wire[15:0] addr_remain3_3815;
address_decode_4 decoder_3_3815 = address_decode_4(addr_selector2_238[7],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3815,addr_remain3_3815);


wire[15:0] addr_selector3_3816;
wire[15:0] addr_remain3_3816;
address_decode_4 decoder_3_3816 = address_decode_4(addr_selector2_238[8],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3816,addr_remain3_3816);


wire[15:0] addr_selector3_3817;
wire[15:0] addr_remain3_3817;
address_decode_4 decoder_3_3817 = address_decode_4(addr_selector2_238[9],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3817,addr_remain3_3817);


wire[15:0] addr_selector3_3818;
wire[15:0] addr_remain3_3818;
address_decode_4 decoder_3_3818 = address_decode_4(addr_selector2_238[10],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3818,addr_remain3_3818);


wire[15:0] addr_selector3_3819;
wire[15:0] addr_remain3_3819;
address_decode_4 decoder_3_3819 = address_decode_4(addr_selector2_238[11],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3819,addr_remain3_3819);


wire[15:0] addr_selector3_3820;
wire[15:0] addr_remain3_3820;
address_decode_4 decoder_3_3820 = address_decode_4(addr_selector2_238[12],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3820,addr_remain3_3820);


wire[15:0] addr_selector3_3821;
wire[15:0] addr_remain3_3821;
address_decode_4 decoder_3_3821 = address_decode_4(addr_selector2_238[13],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3821,addr_remain3_3821);


wire[15:0] addr_selector3_3822;
wire[15:0] addr_remain3_3822;
address_decode_4 decoder_3_3822 = address_decode_4(addr_selector2_238[14],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3822,addr_remain3_3822);


wire[15:0] addr_selector3_3823;
wire[15:0] addr_remain3_3823;
address_decode_4 decoder_3_3823 = address_decode_4(addr_selector2_238[15],addr_remain2_238[15:0],addr_remain2_238,addr_selector3_3823,addr_remain3_3823);


wire[15:0] addr_selector3_3824;
wire[15:0] addr_remain3_3824;
address_decode_4 decoder_3_3824 = address_decode_4(addr_selector2_239[0],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3824,addr_remain3_3824);


wire[15:0] addr_selector3_3825;
wire[15:0] addr_remain3_3825;
address_decode_4 decoder_3_3825 = address_decode_4(addr_selector2_239[1],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3825,addr_remain3_3825);


wire[15:0] addr_selector3_3826;
wire[15:0] addr_remain3_3826;
address_decode_4 decoder_3_3826 = address_decode_4(addr_selector2_239[2],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3826,addr_remain3_3826);


wire[15:0] addr_selector3_3827;
wire[15:0] addr_remain3_3827;
address_decode_4 decoder_3_3827 = address_decode_4(addr_selector2_239[3],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3827,addr_remain3_3827);


wire[15:0] addr_selector3_3828;
wire[15:0] addr_remain3_3828;
address_decode_4 decoder_3_3828 = address_decode_4(addr_selector2_239[4],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3828,addr_remain3_3828);


wire[15:0] addr_selector3_3829;
wire[15:0] addr_remain3_3829;
address_decode_4 decoder_3_3829 = address_decode_4(addr_selector2_239[5],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3829,addr_remain3_3829);


wire[15:0] addr_selector3_3830;
wire[15:0] addr_remain3_3830;
address_decode_4 decoder_3_3830 = address_decode_4(addr_selector2_239[6],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3830,addr_remain3_3830);


wire[15:0] addr_selector3_3831;
wire[15:0] addr_remain3_3831;
address_decode_4 decoder_3_3831 = address_decode_4(addr_selector2_239[7],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3831,addr_remain3_3831);


wire[15:0] addr_selector3_3832;
wire[15:0] addr_remain3_3832;
address_decode_4 decoder_3_3832 = address_decode_4(addr_selector2_239[8],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3832,addr_remain3_3832);


wire[15:0] addr_selector3_3833;
wire[15:0] addr_remain3_3833;
address_decode_4 decoder_3_3833 = address_decode_4(addr_selector2_239[9],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3833,addr_remain3_3833);


wire[15:0] addr_selector3_3834;
wire[15:0] addr_remain3_3834;
address_decode_4 decoder_3_3834 = address_decode_4(addr_selector2_239[10],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3834,addr_remain3_3834);


wire[15:0] addr_selector3_3835;
wire[15:0] addr_remain3_3835;
address_decode_4 decoder_3_3835 = address_decode_4(addr_selector2_239[11],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3835,addr_remain3_3835);


wire[15:0] addr_selector3_3836;
wire[15:0] addr_remain3_3836;
address_decode_4 decoder_3_3836 = address_decode_4(addr_selector2_239[12],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3836,addr_remain3_3836);


wire[15:0] addr_selector3_3837;
wire[15:0] addr_remain3_3837;
address_decode_4 decoder_3_3837 = address_decode_4(addr_selector2_239[13],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3837,addr_remain3_3837);


wire[15:0] addr_selector3_3838;
wire[15:0] addr_remain3_3838;
address_decode_4 decoder_3_3838 = address_decode_4(addr_selector2_239[14],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3838,addr_remain3_3838);


wire[15:0] addr_selector3_3839;
wire[15:0] addr_remain3_3839;
address_decode_4 decoder_3_3839 = address_decode_4(addr_selector2_239[15],addr_remain2_239[15:0],addr_remain2_239,addr_selector3_3839,addr_remain3_3839);


wire[15:0] addr_selector3_3840;
wire[15:0] addr_remain3_3840;
address_decode_4 decoder_3_3840 = address_decode_4(addr_selector2_240[0],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3840,addr_remain3_3840);


wire[15:0] addr_selector3_3841;
wire[15:0] addr_remain3_3841;
address_decode_4 decoder_3_3841 = address_decode_4(addr_selector2_240[1],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3841,addr_remain3_3841);


wire[15:0] addr_selector3_3842;
wire[15:0] addr_remain3_3842;
address_decode_4 decoder_3_3842 = address_decode_4(addr_selector2_240[2],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3842,addr_remain3_3842);


wire[15:0] addr_selector3_3843;
wire[15:0] addr_remain3_3843;
address_decode_4 decoder_3_3843 = address_decode_4(addr_selector2_240[3],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3843,addr_remain3_3843);


wire[15:0] addr_selector3_3844;
wire[15:0] addr_remain3_3844;
address_decode_4 decoder_3_3844 = address_decode_4(addr_selector2_240[4],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3844,addr_remain3_3844);


wire[15:0] addr_selector3_3845;
wire[15:0] addr_remain3_3845;
address_decode_4 decoder_3_3845 = address_decode_4(addr_selector2_240[5],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3845,addr_remain3_3845);


wire[15:0] addr_selector3_3846;
wire[15:0] addr_remain3_3846;
address_decode_4 decoder_3_3846 = address_decode_4(addr_selector2_240[6],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3846,addr_remain3_3846);


wire[15:0] addr_selector3_3847;
wire[15:0] addr_remain3_3847;
address_decode_4 decoder_3_3847 = address_decode_4(addr_selector2_240[7],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3847,addr_remain3_3847);


wire[15:0] addr_selector3_3848;
wire[15:0] addr_remain3_3848;
address_decode_4 decoder_3_3848 = address_decode_4(addr_selector2_240[8],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3848,addr_remain3_3848);


wire[15:0] addr_selector3_3849;
wire[15:0] addr_remain3_3849;
address_decode_4 decoder_3_3849 = address_decode_4(addr_selector2_240[9],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3849,addr_remain3_3849);


wire[15:0] addr_selector3_3850;
wire[15:0] addr_remain3_3850;
address_decode_4 decoder_3_3850 = address_decode_4(addr_selector2_240[10],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3850,addr_remain3_3850);


wire[15:0] addr_selector3_3851;
wire[15:0] addr_remain3_3851;
address_decode_4 decoder_3_3851 = address_decode_4(addr_selector2_240[11],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3851,addr_remain3_3851);


wire[15:0] addr_selector3_3852;
wire[15:0] addr_remain3_3852;
address_decode_4 decoder_3_3852 = address_decode_4(addr_selector2_240[12],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3852,addr_remain3_3852);


wire[15:0] addr_selector3_3853;
wire[15:0] addr_remain3_3853;
address_decode_4 decoder_3_3853 = address_decode_4(addr_selector2_240[13],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3853,addr_remain3_3853);


wire[15:0] addr_selector3_3854;
wire[15:0] addr_remain3_3854;
address_decode_4 decoder_3_3854 = address_decode_4(addr_selector2_240[14],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3854,addr_remain3_3854);


wire[15:0] addr_selector3_3855;
wire[15:0] addr_remain3_3855;
address_decode_4 decoder_3_3855 = address_decode_4(addr_selector2_240[15],addr_remain2_240[15:0],addr_remain2_240,addr_selector3_3855,addr_remain3_3855);


wire[15:0] addr_selector3_3856;
wire[15:0] addr_remain3_3856;
address_decode_4 decoder_3_3856 = address_decode_4(addr_selector2_241[0],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3856,addr_remain3_3856);


wire[15:0] addr_selector3_3857;
wire[15:0] addr_remain3_3857;
address_decode_4 decoder_3_3857 = address_decode_4(addr_selector2_241[1],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3857,addr_remain3_3857);


wire[15:0] addr_selector3_3858;
wire[15:0] addr_remain3_3858;
address_decode_4 decoder_3_3858 = address_decode_4(addr_selector2_241[2],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3858,addr_remain3_3858);


wire[15:0] addr_selector3_3859;
wire[15:0] addr_remain3_3859;
address_decode_4 decoder_3_3859 = address_decode_4(addr_selector2_241[3],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3859,addr_remain3_3859);


wire[15:0] addr_selector3_3860;
wire[15:0] addr_remain3_3860;
address_decode_4 decoder_3_3860 = address_decode_4(addr_selector2_241[4],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3860,addr_remain3_3860);


wire[15:0] addr_selector3_3861;
wire[15:0] addr_remain3_3861;
address_decode_4 decoder_3_3861 = address_decode_4(addr_selector2_241[5],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3861,addr_remain3_3861);


wire[15:0] addr_selector3_3862;
wire[15:0] addr_remain3_3862;
address_decode_4 decoder_3_3862 = address_decode_4(addr_selector2_241[6],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3862,addr_remain3_3862);


wire[15:0] addr_selector3_3863;
wire[15:0] addr_remain3_3863;
address_decode_4 decoder_3_3863 = address_decode_4(addr_selector2_241[7],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3863,addr_remain3_3863);


wire[15:0] addr_selector3_3864;
wire[15:0] addr_remain3_3864;
address_decode_4 decoder_3_3864 = address_decode_4(addr_selector2_241[8],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3864,addr_remain3_3864);


wire[15:0] addr_selector3_3865;
wire[15:0] addr_remain3_3865;
address_decode_4 decoder_3_3865 = address_decode_4(addr_selector2_241[9],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3865,addr_remain3_3865);


wire[15:0] addr_selector3_3866;
wire[15:0] addr_remain3_3866;
address_decode_4 decoder_3_3866 = address_decode_4(addr_selector2_241[10],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3866,addr_remain3_3866);


wire[15:0] addr_selector3_3867;
wire[15:0] addr_remain3_3867;
address_decode_4 decoder_3_3867 = address_decode_4(addr_selector2_241[11],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3867,addr_remain3_3867);


wire[15:0] addr_selector3_3868;
wire[15:0] addr_remain3_3868;
address_decode_4 decoder_3_3868 = address_decode_4(addr_selector2_241[12],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3868,addr_remain3_3868);


wire[15:0] addr_selector3_3869;
wire[15:0] addr_remain3_3869;
address_decode_4 decoder_3_3869 = address_decode_4(addr_selector2_241[13],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3869,addr_remain3_3869);


wire[15:0] addr_selector3_3870;
wire[15:0] addr_remain3_3870;
address_decode_4 decoder_3_3870 = address_decode_4(addr_selector2_241[14],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3870,addr_remain3_3870);


wire[15:0] addr_selector3_3871;
wire[15:0] addr_remain3_3871;
address_decode_4 decoder_3_3871 = address_decode_4(addr_selector2_241[15],addr_remain2_241[15:0],addr_remain2_241,addr_selector3_3871,addr_remain3_3871);


wire[15:0] addr_selector3_3872;
wire[15:0] addr_remain3_3872;
address_decode_4 decoder_3_3872 = address_decode_4(addr_selector2_242[0],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3872,addr_remain3_3872);


wire[15:0] addr_selector3_3873;
wire[15:0] addr_remain3_3873;
address_decode_4 decoder_3_3873 = address_decode_4(addr_selector2_242[1],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3873,addr_remain3_3873);


wire[15:0] addr_selector3_3874;
wire[15:0] addr_remain3_3874;
address_decode_4 decoder_3_3874 = address_decode_4(addr_selector2_242[2],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3874,addr_remain3_3874);


wire[15:0] addr_selector3_3875;
wire[15:0] addr_remain3_3875;
address_decode_4 decoder_3_3875 = address_decode_4(addr_selector2_242[3],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3875,addr_remain3_3875);


wire[15:0] addr_selector3_3876;
wire[15:0] addr_remain3_3876;
address_decode_4 decoder_3_3876 = address_decode_4(addr_selector2_242[4],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3876,addr_remain3_3876);


wire[15:0] addr_selector3_3877;
wire[15:0] addr_remain3_3877;
address_decode_4 decoder_3_3877 = address_decode_4(addr_selector2_242[5],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3877,addr_remain3_3877);


wire[15:0] addr_selector3_3878;
wire[15:0] addr_remain3_3878;
address_decode_4 decoder_3_3878 = address_decode_4(addr_selector2_242[6],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3878,addr_remain3_3878);


wire[15:0] addr_selector3_3879;
wire[15:0] addr_remain3_3879;
address_decode_4 decoder_3_3879 = address_decode_4(addr_selector2_242[7],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3879,addr_remain3_3879);


wire[15:0] addr_selector3_3880;
wire[15:0] addr_remain3_3880;
address_decode_4 decoder_3_3880 = address_decode_4(addr_selector2_242[8],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3880,addr_remain3_3880);


wire[15:0] addr_selector3_3881;
wire[15:0] addr_remain3_3881;
address_decode_4 decoder_3_3881 = address_decode_4(addr_selector2_242[9],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3881,addr_remain3_3881);


wire[15:0] addr_selector3_3882;
wire[15:0] addr_remain3_3882;
address_decode_4 decoder_3_3882 = address_decode_4(addr_selector2_242[10],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3882,addr_remain3_3882);


wire[15:0] addr_selector3_3883;
wire[15:0] addr_remain3_3883;
address_decode_4 decoder_3_3883 = address_decode_4(addr_selector2_242[11],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3883,addr_remain3_3883);


wire[15:0] addr_selector3_3884;
wire[15:0] addr_remain3_3884;
address_decode_4 decoder_3_3884 = address_decode_4(addr_selector2_242[12],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3884,addr_remain3_3884);


wire[15:0] addr_selector3_3885;
wire[15:0] addr_remain3_3885;
address_decode_4 decoder_3_3885 = address_decode_4(addr_selector2_242[13],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3885,addr_remain3_3885);


wire[15:0] addr_selector3_3886;
wire[15:0] addr_remain3_3886;
address_decode_4 decoder_3_3886 = address_decode_4(addr_selector2_242[14],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3886,addr_remain3_3886);


wire[15:0] addr_selector3_3887;
wire[15:0] addr_remain3_3887;
address_decode_4 decoder_3_3887 = address_decode_4(addr_selector2_242[15],addr_remain2_242[15:0],addr_remain2_242,addr_selector3_3887,addr_remain3_3887);


wire[15:0] addr_selector3_3888;
wire[15:0] addr_remain3_3888;
address_decode_4 decoder_3_3888 = address_decode_4(addr_selector2_243[0],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3888,addr_remain3_3888);


wire[15:0] addr_selector3_3889;
wire[15:0] addr_remain3_3889;
address_decode_4 decoder_3_3889 = address_decode_4(addr_selector2_243[1],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3889,addr_remain3_3889);


wire[15:0] addr_selector3_3890;
wire[15:0] addr_remain3_3890;
address_decode_4 decoder_3_3890 = address_decode_4(addr_selector2_243[2],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3890,addr_remain3_3890);


wire[15:0] addr_selector3_3891;
wire[15:0] addr_remain3_3891;
address_decode_4 decoder_3_3891 = address_decode_4(addr_selector2_243[3],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3891,addr_remain3_3891);


wire[15:0] addr_selector3_3892;
wire[15:0] addr_remain3_3892;
address_decode_4 decoder_3_3892 = address_decode_4(addr_selector2_243[4],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3892,addr_remain3_3892);


wire[15:0] addr_selector3_3893;
wire[15:0] addr_remain3_3893;
address_decode_4 decoder_3_3893 = address_decode_4(addr_selector2_243[5],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3893,addr_remain3_3893);


wire[15:0] addr_selector3_3894;
wire[15:0] addr_remain3_3894;
address_decode_4 decoder_3_3894 = address_decode_4(addr_selector2_243[6],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3894,addr_remain3_3894);


wire[15:0] addr_selector3_3895;
wire[15:0] addr_remain3_3895;
address_decode_4 decoder_3_3895 = address_decode_4(addr_selector2_243[7],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3895,addr_remain3_3895);


wire[15:0] addr_selector3_3896;
wire[15:0] addr_remain3_3896;
address_decode_4 decoder_3_3896 = address_decode_4(addr_selector2_243[8],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3896,addr_remain3_3896);


wire[15:0] addr_selector3_3897;
wire[15:0] addr_remain3_3897;
address_decode_4 decoder_3_3897 = address_decode_4(addr_selector2_243[9],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3897,addr_remain3_3897);


wire[15:0] addr_selector3_3898;
wire[15:0] addr_remain3_3898;
address_decode_4 decoder_3_3898 = address_decode_4(addr_selector2_243[10],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3898,addr_remain3_3898);


wire[15:0] addr_selector3_3899;
wire[15:0] addr_remain3_3899;
address_decode_4 decoder_3_3899 = address_decode_4(addr_selector2_243[11],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3899,addr_remain3_3899);


wire[15:0] addr_selector3_3900;
wire[15:0] addr_remain3_3900;
address_decode_4 decoder_3_3900 = address_decode_4(addr_selector2_243[12],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3900,addr_remain3_3900);


wire[15:0] addr_selector3_3901;
wire[15:0] addr_remain3_3901;
address_decode_4 decoder_3_3901 = address_decode_4(addr_selector2_243[13],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3901,addr_remain3_3901);


wire[15:0] addr_selector3_3902;
wire[15:0] addr_remain3_3902;
address_decode_4 decoder_3_3902 = address_decode_4(addr_selector2_243[14],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3902,addr_remain3_3902);


wire[15:0] addr_selector3_3903;
wire[15:0] addr_remain3_3903;
address_decode_4 decoder_3_3903 = address_decode_4(addr_selector2_243[15],addr_remain2_243[15:0],addr_remain2_243,addr_selector3_3903,addr_remain3_3903);


wire[15:0] addr_selector3_3904;
wire[15:0] addr_remain3_3904;
address_decode_4 decoder_3_3904 = address_decode_4(addr_selector2_244[0],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3904,addr_remain3_3904);


wire[15:0] addr_selector3_3905;
wire[15:0] addr_remain3_3905;
address_decode_4 decoder_3_3905 = address_decode_4(addr_selector2_244[1],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3905,addr_remain3_3905);


wire[15:0] addr_selector3_3906;
wire[15:0] addr_remain3_3906;
address_decode_4 decoder_3_3906 = address_decode_4(addr_selector2_244[2],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3906,addr_remain3_3906);


wire[15:0] addr_selector3_3907;
wire[15:0] addr_remain3_3907;
address_decode_4 decoder_3_3907 = address_decode_4(addr_selector2_244[3],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3907,addr_remain3_3907);


wire[15:0] addr_selector3_3908;
wire[15:0] addr_remain3_3908;
address_decode_4 decoder_3_3908 = address_decode_4(addr_selector2_244[4],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3908,addr_remain3_3908);


wire[15:0] addr_selector3_3909;
wire[15:0] addr_remain3_3909;
address_decode_4 decoder_3_3909 = address_decode_4(addr_selector2_244[5],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3909,addr_remain3_3909);


wire[15:0] addr_selector3_3910;
wire[15:0] addr_remain3_3910;
address_decode_4 decoder_3_3910 = address_decode_4(addr_selector2_244[6],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3910,addr_remain3_3910);


wire[15:0] addr_selector3_3911;
wire[15:0] addr_remain3_3911;
address_decode_4 decoder_3_3911 = address_decode_4(addr_selector2_244[7],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3911,addr_remain3_3911);


wire[15:0] addr_selector3_3912;
wire[15:0] addr_remain3_3912;
address_decode_4 decoder_3_3912 = address_decode_4(addr_selector2_244[8],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3912,addr_remain3_3912);


wire[15:0] addr_selector3_3913;
wire[15:0] addr_remain3_3913;
address_decode_4 decoder_3_3913 = address_decode_4(addr_selector2_244[9],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3913,addr_remain3_3913);


wire[15:0] addr_selector3_3914;
wire[15:0] addr_remain3_3914;
address_decode_4 decoder_3_3914 = address_decode_4(addr_selector2_244[10],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3914,addr_remain3_3914);


wire[15:0] addr_selector3_3915;
wire[15:0] addr_remain3_3915;
address_decode_4 decoder_3_3915 = address_decode_4(addr_selector2_244[11],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3915,addr_remain3_3915);


wire[15:0] addr_selector3_3916;
wire[15:0] addr_remain3_3916;
address_decode_4 decoder_3_3916 = address_decode_4(addr_selector2_244[12],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3916,addr_remain3_3916);


wire[15:0] addr_selector3_3917;
wire[15:0] addr_remain3_3917;
address_decode_4 decoder_3_3917 = address_decode_4(addr_selector2_244[13],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3917,addr_remain3_3917);


wire[15:0] addr_selector3_3918;
wire[15:0] addr_remain3_3918;
address_decode_4 decoder_3_3918 = address_decode_4(addr_selector2_244[14],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3918,addr_remain3_3918);


wire[15:0] addr_selector3_3919;
wire[15:0] addr_remain3_3919;
address_decode_4 decoder_3_3919 = address_decode_4(addr_selector2_244[15],addr_remain2_244[15:0],addr_remain2_244,addr_selector3_3919,addr_remain3_3919);


wire[15:0] addr_selector3_3920;
wire[15:0] addr_remain3_3920;
address_decode_4 decoder_3_3920 = address_decode_4(addr_selector2_245[0],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3920,addr_remain3_3920);


wire[15:0] addr_selector3_3921;
wire[15:0] addr_remain3_3921;
address_decode_4 decoder_3_3921 = address_decode_4(addr_selector2_245[1],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3921,addr_remain3_3921);


wire[15:0] addr_selector3_3922;
wire[15:0] addr_remain3_3922;
address_decode_4 decoder_3_3922 = address_decode_4(addr_selector2_245[2],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3922,addr_remain3_3922);


wire[15:0] addr_selector3_3923;
wire[15:0] addr_remain3_3923;
address_decode_4 decoder_3_3923 = address_decode_4(addr_selector2_245[3],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3923,addr_remain3_3923);


wire[15:0] addr_selector3_3924;
wire[15:0] addr_remain3_3924;
address_decode_4 decoder_3_3924 = address_decode_4(addr_selector2_245[4],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3924,addr_remain3_3924);


wire[15:0] addr_selector3_3925;
wire[15:0] addr_remain3_3925;
address_decode_4 decoder_3_3925 = address_decode_4(addr_selector2_245[5],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3925,addr_remain3_3925);


wire[15:0] addr_selector3_3926;
wire[15:0] addr_remain3_3926;
address_decode_4 decoder_3_3926 = address_decode_4(addr_selector2_245[6],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3926,addr_remain3_3926);


wire[15:0] addr_selector3_3927;
wire[15:0] addr_remain3_3927;
address_decode_4 decoder_3_3927 = address_decode_4(addr_selector2_245[7],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3927,addr_remain3_3927);


wire[15:0] addr_selector3_3928;
wire[15:0] addr_remain3_3928;
address_decode_4 decoder_3_3928 = address_decode_4(addr_selector2_245[8],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3928,addr_remain3_3928);


wire[15:0] addr_selector3_3929;
wire[15:0] addr_remain3_3929;
address_decode_4 decoder_3_3929 = address_decode_4(addr_selector2_245[9],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3929,addr_remain3_3929);


wire[15:0] addr_selector3_3930;
wire[15:0] addr_remain3_3930;
address_decode_4 decoder_3_3930 = address_decode_4(addr_selector2_245[10],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3930,addr_remain3_3930);


wire[15:0] addr_selector3_3931;
wire[15:0] addr_remain3_3931;
address_decode_4 decoder_3_3931 = address_decode_4(addr_selector2_245[11],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3931,addr_remain3_3931);


wire[15:0] addr_selector3_3932;
wire[15:0] addr_remain3_3932;
address_decode_4 decoder_3_3932 = address_decode_4(addr_selector2_245[12],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3932,addr_remain3_3932);


wire[15:0] addr_selector3_3933;
wire[15:0] addr_remain3_3933;
address_decode_4 decoder_3_3933 = address_decode_4(addr_selector2_245[13],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3933,addr_remain3_3933);


wire[15:0] addr_selector3_3934;
wire[15:0] addr_remain3_3934;
address_decode_4 decoder_3_3934 = address_decode_4(addr_selector2_245[14],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3934,addr_remain3_3934);


wire[15:0] addr_selector3_3935;
wire[15:0] addr_remain3_3935;
address_decode_4 decoder_3_3935 = address_decode_4(addr_selector2_245[15],addr_remain2_245[15:0],addr_remain2_245,addr_selector3_3935,addr_remain3_3935);


wire[15:0] addr_selector3_3936;
wire[15:0] addr_remain3_3936;
address_decode_4 decoder_3_3936 = address_decode_4(addr_selector2_246[0],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3936,addr_remain3_3936);


wire[15:0] addr_selector3_3937;
wire[15:0] addr_remain3_3937;
address_decode_4 decoder_3_3937 = address_decode_4(addr_selector2_246[1],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3937,addr_remain3_3937);


wire[15:0] addr_selector3_3938;
wire[15:0] addr_remain3_3938;
address_decode_4 decoder_3_3938 = address_decode_4(addr_selector2_246[2],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3938,addr_remain3_3938);


wire[15:0] addr_selector3_3939;
wire[15:0] addr_remain3_3939;
address_decode_4 decoder_3_3939 = address_decode_4(addr_selector2_246[3],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3939,addr_remain3_3939);


wire[15:0] addr_selector3_3940;
wire[15:0] addr_remain3_3940;
address_decode_4 decoder_3_3940 = address_decode_4(addr_selector2_246[4],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3940,addr_remain3_3940);


wire[15:0] addr_selector3_3941;
wire[15:0] addr_remain3_3941;
address_decode_4 decoder_3_3941 = address_decode_4(addr_selector2_246[5],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3941,addr_remain3_3941);


wire[15:0] addr_selector3_3942;
wire[15:0] addr_remain3_3942;
address_decode_4 decoder_3_3942 = address_decode_4(addr_selector2_246[6],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3942,addr_remain3_3942);


wire[15:0] addr_selector3_3943;
wire[15:0] addr_remain3_3943;
address_decode_4 decoder_3_3943 = address_decode_4(addr_selector2_246[7],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3943,addr_remain3_3943);


wire[15:0] addr_selector3_3944;
wire[15:0] addr_remain3_3944;
address_decode_4 decoder_3_3944 = address_decode_4(addr_selector2_246[8],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3944,addr_remain3_3944);


wire[15:0] addr_selector3_3945;
wire[15:0] addr_remain3_3945;
address_decode_4 decoder_3_3945 = address_decode_4(addr_selector2_246[9],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3945,addr_remain3_3945);


wire[15:0] addr_selector3_3946;
wire[15:0] addr_remain3_3946;
address_decode_4 decoder_3_3946 = address_decode_4(addr_selector2_246[10],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3946,addr_remain3_3946);


wire[15:0] addr_selector3_3947;
wire[15:0] addr_remain3_3947;
address_decode_4 decoder_3_3947 = address_decode_4(addr_selector2_246[11],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3947,addr_remain3_3947);


wire[15:0] addr_selector3_3948;
wire[15:0] addr_remain3_3948;
address_decode_4 decoder_3_3948 = address_decode_4(addr_selector2_246[12],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3948,addr_remain3_3948);


wire[15:0] addr_selector3_3949;
wire[15:0] addr_remain3_3949;
address_decode_4 decoder_3_3949 = address_decode_4(addr_selector2_246[13],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3949,addr_remain3_3949);


wire[15:0] addr_selector3_3950;
wire[15:0] addr_remain3_3950;
address_decode_4 decoder_3_3950 = address_decode_4(addr_selector2_246[14],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3950,addr_remain3_3950);


wire[15:0] addr_selector3_3951;
wire[15:0] addr_remain3_3951;
address_decode_4 decoder_3_3951 = address_decode_4(addr_selector2_246[15],addr_remain2_246[15:0],addr_remain2_246,addr_selector3_3951,addr_remain3_3951);


wire[15:0] addr_selector3_3952;
wire[15:0] addr_remain3_3952;
address_decode_4 decoder_3_3952 = address_decode_4(addr_selector2_247[0],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3952,addr_remain3_3952);


wire[15:0] addr_selector3_3953;
wire[15:0] addr_remain3_3953;
address_decode_4 decoder_3_3953 = address_decode_4(addr_selector2_247[1],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3953,addr_remain3_3953);


wire[15:0] addr_selector3_3954;
wire[15:0] addr_remain3_3954;
address_decode_4 decoder_3_3954 = address_decode_4(addr_selector2_247[2],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3954,addr_remain3_3954);


wire[15:0] addr_selector3_3955;
wire[15:0] addr_remain3_3955;
address_decode_4 decoder_3_3955 = address_decode_4(addr_selector2_247[3],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3955,addr_remain3_3955);


wire[15:0] addr_selector3_3956;
wire[15:0] addr_remain3_3956;
address_decode_4 decoder_3_3956 = address_decode_4(addr_selector2_247[4],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3956,addr_remain3_3956);


wire[15:0] addr_selector3_3957;
wire[15:0] addr_remain3_3957;
address_decode_4 decoder_3_3957 = address_decode_4(addr_selector2_247[5],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3957,addr_remain3_3957);


wire[15:0] addr_selector3_3958;
wire[15:0] addr_remain3_3958;
address_decode_4 decoder_3_3958 = address_decode_4(addr_selector2_247[6],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3958,addr_remain3_3958);


wire[15:0] addr_selector3_3959;
wire[15:0] addr_remain3_3959;
address_decode_4 decoder_3_3959 = address_decode_4(addr_selector2_247[7],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3959,addr_remain3_3959);


wire[15:0] addr_selector3_3960;
wire[15:0] addr_remain3_3960;
address_decode_4 decoder_3_3960 = address_decode_4(addr_selector2_247[8],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3960,addr_remain3_3960);


wire[15:0] addr_selector3_3961;
wire[15:0] addr_remain3_3961;
address_decode_4 decoder_3_3961 = address_decode_4(addr_selector2_247[9],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3961,addr_remain3_3961);


wire[15:0] addr_selector3_3962;
wire[15:0] addr_remain3_3962;
address_decode_4 decoder_3_3962 = address_decode_4(addr_selector2_247[10],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3962,addr_remain3_3962);


wire[15:0] addr_selector3_3963;
wire[15:0] addr_remain3_3963;
address_decode_4 decoder_3_3963 = address_decode_4(addr_selector2_247[11],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3963,addr_remain3_3963);


wire[15:0] addr_selector3_3964;
wire[15:0] addr_remain3_3964;
address_decode_4 decoder_3_3964 = address_decode_4(addr_selector2_247[12],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3964,addr_remain3_3964);


wire[15:0] addr_selector3_3965;
wire[15:0] addr_remain3_3965;
address_decode_4 decoder_3_3965 = address_decode_4(addr_selector2_247[13],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3965,addr_remain3_3965);


wire[15:0] addr_selector3_3966;
wire[15:0] addr_remain3_3966;
address_decode_4 decoder_3_3966 = address_decode_4(addr_selector2_247[14],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3966,addr_remain3_3966);


wire[15:0] addr_selector3_3967;
wire[15:0] addr_remain3_3967;
address_decode_4 decoder_3_3967 = address_decode_4(addr_selector2_247[15],addr_remain2_247[15:0],addr_remain2_247,addr_selector3_3967,addr_remain3_3967);


wire[15:0] addr_selector3_3968;
wire[15:0] addr_remain3_3968;
address_decode_4 decoder_3_3968 = address_decode_4(addr_selector2_248[0],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3968,addr_remain3_3968);


wire[15:0] addr_selector3_3969;
wire[15:0] addr_remain3_3969;
address_decode_4 decoder_3_3969 = address_decode_4(addr_selector2_248[1],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3969,addr_remain3_3969);


wire[15:0] addr_selector3_3970;
wire[15:0] addr_remain3_3970;
address_decode_4 decoder_3_3970 = address_decode_4(addr_selector2_248[2],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3970,addr_remain3_3970);


wire[15:0] addr_selector3_3971;
wire[15:0] addr_remain3_3971;
address_decode_4 decoder_3_3971 = address_decode_4(addr_selector2_248[3],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3971,addr_remain3_3971);


wire[15:0] addr_selector3_3972;
wire[15:0] addr_remain3_3972;
address_decode_4 decoder_3_3972 = address_decode_4(addr_selector2_248[4],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3972,addr_remain3_3972);


wire[15:0] addr_selector3_3973;
wire[15:0] addr_remain3_3973;
address_decode_4 decoder_3_3973 = address_decode_4(addr_selector2_248[5],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3973,addr_remain3_3973);


wire[15:0] addr_selector3_3974;
wire[15:0] addr_remain3_3974;
address_decode_4 decoder_3_3974 = address_decode_4(addr_selector2_248[6],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3974,addr_remain3_3974);


wire[15:0] addr_selector3_3975;
wire[15:0] addr_remain3_3975;
address_decode_4 decoder_3_3975 = address_decode_4(addr_selector2_248[7],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3975,addr_remain3_3975);


wire[15:0] addr_selector3_3976;
wire[15:0] addr_remain3_3976;
address_decode_4 decoder_3_3976 = address_decode_4(addr_selector2_248[8],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3976,addr_remain3_3976);


wire[15:0] addr_selector3_3977;
wire[15:0] addr_remain3_3977;
address_decode_4 decoder_3_3977 = address_decode_4(addr_selector2_248[9],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3977,addr_remain3_3977);


wire[15:0] addr_selector3_3978;
wire[15:0] addr_remain3_3978;
address_decode_4 decoder_3_3978 = address_decode_4(addr_selector2_248[10],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3978,addr_remain3_3978);


wire[15:0] addr_selector3_3979;
wire[15:0] addr_remain3_3979;
address_decode_4 decoder_3_3979 = address_decode_4(addr_selector2_248[11],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3979,addr_remain3_3979);


wire[15:0] addr_selector3_3980;
wire[15:0] addr_remain3_3980;
address_decode_4 decoder_3_3980 = address_decode_4(addr_selector2_248[12],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3980,addr_remain3_3980);


wire[15:0] addr_selector3_3981;
wire[15:0] addr_remain3_3981;
address_decode_4 decoder_3_3981 = address_decode_4(addr_selector2_248[13],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3981,addr_remain3_3981);


wire[15:0] addr_selector3_3982;
wire[15:0] addr_remain3_3982;
address_decode_4 decoder_3_3982 = address_decode_4(addr_selector2_248[14],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3982,addr_remain3_3982);


wire[15:0] addr_selector3_3983;
wire[15:0] addr_remain3_3983;
address_decode_4 decoder_3_3983 = address_decode_4(addr_selector2_248[15],addr_remain2_248[15:0],addr_remain2_248,addr_selector3_3983,addr_remain3_3983);


wire[15:0] addr_selector3_3984;
wire[15:0] addr_remain3_3984;
address_decode_4 decoder_3_3984 = address_decode_4(addr_selector2_249[0],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3984,addr_remain3_3984);


wire[15:0] addr_selector3_3985;
wire[15:0] addr_remain3_3985;
address_decode_4 decoder_3_3985 = address_decode_4(addr_selector2_249[1],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3985,addr_remain3_3985);


wire[15:0] addr_selector3_3986;
wire[15:0] addr_remain3_3986;
address_decode_4 decoder_3_3986 = address_decode_4(addr_selector2_249[2],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3986,addr_remain3_3986);


wire[15:0] addr_selector3_3987;
wire[15:0] addr_remain3_3987;
address_decode_4 decoder_3_3987 = address_decode_4(addr_selector2_249[3],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3987,addr_remain3_3987);


wire[15:0] addr_selector3_3988;
wire[15:0] addr_remain3_3988;
address_decode_4 decoder_3_3988 = address_decode_4(addr_selector2_249[4],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3988,addr_remain3_3988);


wire[15:0] addr_selector3_3989;
wire[15:0] addr_remain3_3989;
address_decode_4 decoder_3_3989 = address_decode_4(addr_selector2_249[5],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3989,addr_remain3_3989);


wire[15:0] addr_selector3_3990;
wire[15:0] addr_remain3_3990;
address_decode_4 decoder_3_3990 = address_decode_4(addr_selector2_249[6],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3990,addr_remain3_3990);


wire[15:0] addr_selector3_3991;
wire[15:0] addr_remain3_3991;
address_decode_4 decoder_3_3991 = address_decode_4(addr_selector2_249[7],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3991,addr_remain3_3991);


wire[15:0] addr_selector3_3992;
wire[15:0] addr_remain3_3992;
address_decode_4 decoder_3_3992 = address_decode_4(addr_selector2_249[8],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3992,addr_remain3_3992);


wire[15:0] addr_selector3_3993;
wire[15:0] addr_remain3_3993;
address_decode_4 decoder_3_3993 = address_decode_4(addr_selector2_249[9],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3993,addr_remain3_3993);


wire[15:0] addr_selector3_3994;
wire[15:0] addr_remain3_3994;
address_decode_4 decoder_3_3994 = address_decode_4(addr_selector2_249[10],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3994,addr_remain3_3994);


wire[15:0] addr_selector3_3995;
wire[15:0] addr_remain3_3995;
address_decode_4 decoder_3_3995 = address_decode_4(addr_selector2_249[11],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3995,addr_remain3_3995);


wire[15:0] addr_selector3_3996;
wire[15:0] addr_remain3_3996;
address_decode_4 decoder_3_3996 = address_decode_4(addr_selector2_249[12],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3996,addr_remain3_3996);


wire[15:0] addr_selector3_3997;
wire[15:0] addr_remain3_3997;
address_decode_4 decoder_3_3997 = address_decode_4(addr_selector2_249[13],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3997,addr_remain3_3997);


wire[15:0] addr_selector3_3998;
wire[15:0] addr_remain3_3998;
address_decode_4 decoder_3_3998 = address_decode_4(addr_selector2_249[14],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3998,addr_remain3_3998);


wire[15:0] addr_selector3_3999;
wire[15:0] addr_remain3_3999;
address_decode_4 decoder_3_3999 = address_decode_4(addr_selector2_249[15],addr_remain2_249[15:0],addr_remain2_249,addr_selector3_3999,addr_remain3_3999);


wire[15:0] addr_selector3_4000;
wire[15:0] addr_remain3_4000;
address_decode_4 decoder_3_4000 = address_decode_4(addr_selector2_250[0],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4000,addr_remain3_4000);


wire[15:0] addr_selector3_4001;
wire[15:0] addr_remain3_4001;
address_decode_4 decoder_3_4001 = address_decode_4(addr_selector2_250[1],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4001,addr_remain3_4001);


wire[15:0] addr_selector3_4002;
wire[15:0] addr_remain3_4002;
address_decode_4 decoder_3_4002 = address_decode_4(addr_selector2_250[2],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4002,addr_remain3_4002);


wire[15:0] addr_selector3_4003;
wire[15:0] addr_remain3_4003;
address_decode_4 decoder_3_4003 = address_decode_4(addr_selector2_250[3],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4003,addr_remain3_4003);


wire[15:0] addr_selector3_4004;
wire[15:0] addr_remain3_4004;
address_decode_4 decoder_3_4004 = address_decode_4(addr_selector2_250[4],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4004,addr_remain3_4004);


wire[15:0] addr_selector3_4005;
wire[15:0] addr_remain3_4005;
address_decode_4 decoder_3_4005 = address_decode_4(addr_selector2_250[5],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4005,addr_remain3_4005);


wire[15:0] addr_selector3_4006;
wire[15:0] addr_remain3_4006;
address_decode_4 decoder_3_4006 = address_decode_4(addr_selector2_250[6],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4006,addr_remain3_4006);


wire[15:0] addr_selector3_4007;
wire[15:0] addr_remain3_4007;
address_decode_4 decoder_3_4007 = address_decode_4(addr_selector2_250[7],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4007,addr_remain3_4007);


wire[15:0] addr_selector3_4008;
wire[15:0] addr_remain3_4008;
address_decode_4 decoder_3_4008 = address_decode_4(addr_selector2_250[8],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4008,addr_remain3_4008);


wire[15:0] addr_selector3_4009;
wire[15:0] addr_remain3_4009;
address_decode_4 decoder_3_4009 = address_decode_4(addr_selector2_250[9],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4009,addr_remain3_4009);


wire[15:0] addr_selector3_4010;
wire[15:0] addr_remain3_4010;
address_decode_4 decoder_3_4010 = address_decode_4(addr_selector2_250[10],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4010,addr_remain3_4010);


wire[15:0] addr_selector3_4011;
wire[15:0] addr_remain3_4011;
address_decode_4 decoder_3_4011 = address_decode_4(addr_selector2_250[11],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4011,addr_remain3_4011);


wire[15:0] addr_selector3_4012;
wire[15:0] addr_remain3_4012;
address_decode_4 decoder_3_4012 = address_decode_4(addr_selector2_250[12],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4012,addr_remain3_4012);


wire[15:0] addr_selector3_4013;
wire[15:0] addr_remain3_4013;
address_decode_4 decoder_3_4013 = address_decode_4(addr_selector2_250[13],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4013,addr_remain3_4013);


wire[15:0] addr_selector3_4014;
wire[15:0] addr_remain3_4014;
address_decode_4 decoder_3_4014 = address_decode_4(addr_selector2_250[14],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4014,addr_remain3_4014);


wire[15:0] addr_selector3_4015;
wire[15:0] addr_remain3_4015;
address_decode_4 decoder_3_4015 = address_decode_4(addr_selector2_250[15],addr_remain2_250[15:0],addr_remain2_250,addr_selector3_4015,addr_remain3_4015);


wire[15:0] addr_selector3_4016;
wire[15:0] addr_remain3_4016;
address_decode_4 decoder_3_4016 = address_decode_4(addr_selector2_251[0],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4016,addr_remain3_4016);


wire[15:0] addr_selector3_4017;
wire[15:0] addr_remain3_4017;
address_decode_4 decoder_3_4017 = address_decode_4(addr_selector2_251[1],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4017,addr_remain3_4017);


wire[15:0] addr_selector3_4018;
wire[15:0] addr_remain3_4018;
address_decode_4 decoder_3_4018 = address_decode_4(addr_selector2_251[2],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4018,addr_remain3_4018);


wire[15:0] addr_selector3_4019;
wire[15:0] addr_remain3_4019;
address_decode_4 decoder_3_4019 = address_decode_4(addr_selector2_251[3],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4019,addr_remain3_4019);


wire[15:0] addr_selector3_4020;
wire[15:0] addr_remain3_4020;
address_decode_4 decoder_3_4020 = address_decode_4(addr_selector2_251[4],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4020,addr_remain3_4020);


wire[15:0] addr_selector3_4021;
wire[15:0] addr_remain3_4021;
address_decode_4 decoder_3_4021 = address_decode_4(addr_selector2_251[5],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4021,addr_remain3_4021);


wire[15:0] addr_selector3_4022;
wire[15:0] addr_remain3_4022;
address_decode_4 decoder_3_4022 = address_decode_4(addr_selector2_251[6],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4022,addr_remain3_4022);


wire[15:0] addr_selector3_4023;
wire[15:0] addr_remain3_4023;
address_decode_4 decoder_3_4023 = address_decode_4(addr_selector2_251[7],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4023,addr_remain3_4023);


wire[15:0] addr_selector3_4024;
wire[15:0] addr_remain3_4024;
address_decode_4 decoder_3_4024 = address_decode_4(addr_selector2_251[8],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4024,addr_remain3_4024);


wire[15:0] addr_selector3_4025;
wire[15:0] addr_remain3_4025;
address_decode_4 decoder_3_4025 = address_decode_4(addr_selector2_251[9],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4025,addr_remain3_4025);


wire[15:0] addr_selector3_4026;
wire[15:0] addr_remain3_4026;
address_decode_4 decoder_3_4026 = address_decode_4(addr_selector2_251[10],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4026,addr_remain3_4026);


wire[15:0] addr_selector3_4027;
wire[15:0] addr_remain3_4027;
address_decode_4 decoder_3_4027 = address_decode_4(addr_selector2_251[11],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4027,addr_remain3_4027);


wire[15:0] addr_selector3_4028;
wire[15:0] addr_remain3_4028;
address_decode_4 decoder_3_4028 = address_decode_4(addr_selector2_251[12],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4028,addr_remain3_4028);


wire[15:0] addr_selector3_4029;
wire[15:0] addr_remain3_4029;
address_decode_4 decoder_3_4029 = address_decode_4(addr_selector2_251[13],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4029,addr_remain3_4029);


wire[15:0] addr_selector3_4030;
wire[15:0] addr_remain3_4030;
address_decode_4 decoder_3_4030 = address_decode_4(addr_selector2_251[14],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4030,addr_remain3_4030);


wire[15:0] addr_selector3_4031;
wire[15:0] addr_remain3_4031;
address_decode_4 decoder_3_4031 = address_decode_4(addr_selector2_251[15],addr_remain2_251[15:0],addr_remain2_251,addr_selector3_4031,addr_remain3_4031);


wire[15:0] addr_selector3_4032;
wire[15:0] addr_remain3_4032;
address_decode_4 decoder_3_4032 = address_decode_4(addr_selector2_252[0],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4032,addr_remain3_4032);


wire[15:0] addr_selector3_4033;
wire[15:0] addr_remain3_4033;
address_decode_4 decoder_3_4033 = address_decode_4(addr_selector2_252[1],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4033,addr_remain3_4033);


wire[15:0] addr_selector3_4034;
wire[15:0] addr_remain3_4034;
address_decode_4 decoder_3_4034 = address_decode_4(addr_selector2_252[2],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4034,addr_remain3_4034);


wire[15:0] addr_selector3_4035;
wire[15:0] addr_remain3_4035;
address_decode_4 decoder_3_4035 = address_decode_4(addr_selector2_252[3],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4035,addr_remain3_4035);


wire[15:0] addr_selector3_4036;
wire[15:0] addr_remain3_4036;
address_decode_4 decoder_3_4036 = address_decode_4(addr_selector2_252[4],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4036,addr_remain3_4036);


wire[15:0] addr_selector3_4037;
wire[15:0] addr_remain3_4037;
address_decode_4 decoder_3_4037 = address_decode_4(addr_selector2_252[5],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4037,addr_remain3_4037);


wire[15:0] addr_selector3_4038;
wire[15:0] addr_remain3_4038;
address_decode_4 decoder_3_4038 = address_decode_4(addr_selector2_252[6],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4038,addr_remain3_4038);


wire[15:0] addr_selector3_4039;
wire[15:0] addr_remain3_4039;
address_decode_4 decoder_3_4039 = address_decode_4(addr_selector2_252[7],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4039,addr_remain3_4039);


wire[15:0] addr_selector3_4040;
wire[15:0] addr_remain3_4040;
address_decode_4 decoder_3_4040 = address_decode_4(addr_selector2_252[8],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4040,addr_remain3_4040);


wire[15:0] addr_selector3_4041;
wire[15:0] addr_remain3_4041;
address_decode_4 decoder_3_4041 = address_decode_4(addr_selector2_252[9],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4041,addr_remain3_4041);


wire[15:0] addr_selector3_4042;
wire[15:0] addr_remain3_4042;
address_decode_4 decoder_3_4042 = address_decode_4(addr_selector2_252[10],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4042,addr_remain3_4042);


wire[15:0] addr_selector3_4043;
wire[15:0] addr_remain3_4043;
address_decode_4 decoder_3_4043 = address_decode_4(addr_selector2_252[11],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4043,addr_remain3_4043);


wire[15:0] addr_selector3_4044;
wire[15:0] addr_remain3_4044;
address_decode_4 decoder_3_4044 = address_decode_4(addr_selector2_252[12],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4044,addr_remain3_4044);


wire[15:0] addr_selector3_4045;
wire[15:0] addr_remain3_4045;
address_decode_4 decoder_3_4045 = address_decode_4(addr_selector2_252[13],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4045,addr_remain3_4045);


wire[15:0] addr_selector3_4046;
wire[15:0] addr_remain3_4046;
address_decode_4 decoder_3_4046 = address_decode_4(addr_selector2_252[14],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4046,addr_remain3_4046);


wire[15:0] addr_selector3_4047;
wire[15:0] addr_remain3_4047;
address_decode_4 decoder_3_4047 = address_decode_4(addr_selector2_252[15],addr_remain2_252[15:0],addr_remain2_252,addr_selector3_4047,addr_remain3_4047);


wire[15:0] addr_selector3_4048;
wire[15:0] addr_remain3_4048;
address_decode_4 decoder_3_4048 = address_decode_4(addr_selector2_253[0],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4048,addr_remain3_4048);


wire[15:0] addr_selector3_4049;
wire[15:0] addr_remain3_4049;
address_decode_4 decoder_3_4049 = address_decode_4(addr_selector2_253[1],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4049,addr_remain3_4049);


wire[15:0] addr_selector3_4050;
wire[15:0] addr_remain3_4050;
address_decode_4 decoder_3_4050 = address_decode_4(addr_selector2_253[2],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4050,addr_remain3_4050);


wire[15:0] addr_selector3_4051;
wire[15:0] addr_remain3_4051;
address_decode_4 decoder_3_4051 = address_decode_4(addr_selector2_253[3],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4051,addr_remain3_4051);


wire[15:0] addr_selector3_4052;
wire[15:0] addr_remain3_4052;
address_decode_4 decoder_3_4052 = address_decode_4(addr_selector2_253[4],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4052,addr_remain3_4052);


wire[15:0] addr_selector3_4053;
wire[15:0] addr_remain3_4053;
address_decode_4 decoder_3_4053 = address_decode_4(addr_selector2_253[5],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4053,addr_remain3_4053);


wire[15:0] addr_selector3_4054;
wire[15:0] addr_remain3_4054;
address_decode_4 decoder_3_4054 = address_decode_4(addr_selector2_253[6],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4054,addr_remain3_4054);


wire[15:0] addr_selector3_4055;
wire[15:0] addr_remain3_4055;
address_decode_4 decoder_3_4055 = address_decode_4(addr_selector2_253[7],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4055,addr_remain3_4055);


wire[15:0] addr_selector3_4056;
wire[15:0] addr_remain3_4056;
address_decode_4 decoder_3_4056 = address_decode_4(addr_selector2_253[8],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4056,addr_remain3_4056);


wire[15:0] addr_selector3_4057;
wire[15:0] addr_remain3_4057;
address_decode_4 decoder_3_4057 = address_decode_4(addr_selector2_253[9],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4057,addr_remain3_4057);


wire[15:0] addr_selector3_4058;
wire[15:0] addr_remain3_4058;
address_decode_4 decoder_3_4058 = address_decode_4(addr_selector2_253[10],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4058,addr_remain3_4058);


wire[15:0] addr_selector3_4059;
wire[15:0] addr_remain3_4059;
address_decode_4 decoder_3_4059 = address_decode_4(addr_selector2_253[11],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4059,addr_remain3_4059);


wire[15:0] addr_selector3_4060;
wire[15:0] addr_remain3_4060;
address_decode_4 decoder_3_4060 = address_decode_4(addr_selector2_253[12],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4060,addr_remain3_4060);


wire[15:0] addr_selector3_4061;
wire[15:0] addr_remain3_4061;
address_decode_4 decoder_3_4061 = address_decode_4(addr_selector2_253[13],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4061,addr_remain3_4061);


wire[15:0] addr_selector3_4062;
wire[15:0] addr_remain3_4062;
address_decode_4 decoder_3_4062 = address_decode_4(addr_selector2_253[14],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4062,addr_remain3_4062);


wire[15:0] addr_selector3_4063;
wire[15:0] addr_remain3_4063;
address_decode_4 decoder_3_4063 = address_decode_4(addr_selector2_253[15],addr_remain2_253[15:0],addr_remain2_253,addr_selector3_4063,addr_remain3_4063);


wire[15:0] addr_selector3_4064;
wire[15:0] addr_remain3_4064;
address_decode_4 decoder_3_4064 = address_decode_4(addr_selector2_254[0],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4064,addr_remain3_4064);


wire[15:0] addr_selector3_4065;
wire[15:0] addr_remain3_4065;
address_decode_4 decoder_3_4065 = address_decode_4(addr_selector2_254[1],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4065,addr_remain3_4065);


wire[15:0] addr_selector3_4066;
wire[15:0] addr_remain3_4066;
address_decode_4 decoder_3_4066 = address_decode_4(addr_selector2_254[2],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4066,addr_remain3_4066);


wire[15:0] addr_selector3_4067;
wire[15:0] addr_remain3_4067;
address_decode_4 decoder_3_4067 = address_decode_4(addr_selector2_254[3],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4067,addr_remain3_4067);


wire[15:0] addr_selector3_4068;
wire[15:0] addr_remain3_4068;
address_decode_4 decoder_3_4068 = address_decode_4(addr_selector2_254[4],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4068,addr_remain3_4068);


wire[15:0] addr_selector3_4069;
wire[15:0] addr_remain3_4069;
address_decode_4 decoder_3_4069 = address_decode_4(addr_selector2_254[5],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4069,addr_remain3_4069);


wire[15:0] addr_selector3_4070;
wire[15:0] addr_remain3_4070;
address_decode_4 decoder_3_4070 = address_decode_4(addr_selector2_254[6],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4070,addr_remain3_4070);


wire[15:0] addr_selector3_4071;
wire[15:0] addr_remain3_4071;
address_decode_4 decoder_3_4071 = address_decode_4(addr_selector2_254[7],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4071,addr_remain3_4071);


wire[15:0] addr_selector3_4072;
wire[15:0] addr_remain3_4072;
address_decode_4 decoder_3_4072 = address_decode_4(addr_selector2_254[8],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4072,addr_remain3_4072);


wire[15:0] addr_selector3_4073;
wire[15:0] addr_remain3_4073;
address_decode_4 decoder_3_4073 = address_decode_4(addr_selector2_254[9],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4073,addr_remain3_4073);


wire[15:0] addr_selector3_4074;
wire[15:0] addr_remain3_4074;
address_decode_4 decoder_3_4074 = address_decode_4(addr_selector2_254[10],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4074,addr_remain3_4074);


wire[15:0] addr_selector3_4075;
wire[15:0] addr_remain3_4075;
address_decode_4 decoder_3_4075 = address_decode_4(addr_selector2_254[11],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4075,addr_remain3_4075);


wire[15:0] addr_selector3_4076;
wire[15:0] addr_remain3_4076;
address_decode_4 decoder_3_4076 = address_decode_4(addr_selector2_254[12],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4076,addr_remain3_4076);


wire[15:0] addr_selector3_4077;
wire[15:0] addr_remain3_4077;
address_decode_4 decoder_3_4077 = address_decode_4(addr_selector2_254[13],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4077,addr_remain3_4077);


wire[15:0] addr_selector3_4078;
wire[15:0] addr_remain3_4078;
address_decode_4 decoder_3_4078 = address_decode_4(addr_selector2_254[14],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4078,addr_remain3_4078);


wire[15:0] addr_selector3_4079;
wire[15:0] addr_remain3_4079;
address_decode_4 decoder_3_4079 = address_decode_4(addr_selector2_254[15],addr_remain2_254[15:0],addr_remain2_254,addr_selector3_4079,addr_remain3_4079);


wire[15:0] addr_selector3_4080;
wire[15:0] addr_remain3_4080;
address_decode_4 decoder_3_4080 = address_decode_4(addr_selector2_255[0],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4080,addr_remain3_4080);


wire[15:0] addr_selector3_4081;
wire[15:0] addr_remain3_4081;
address_decode_4 decoder_3_4081 = address_decode_4(addr_selector2_255[1],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4081,addr_remain3_4081);


wire[15:0] addr_selector3_4082;
wire[15:0] addr_remain3_4082;
address_decode_4 decoder_3_4082 = address_decode_4(addr_selector2_255[2],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4082,addr_remain3_4082);


wire[15:0] addr_selector3_4083;
wire[15:0] addr_remain3_4083;
address_decode_4 decoder_3_4083 = address_decode_4(addr_selector2_255[3],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4083,addr_remain3_4083);


wire[15:0] addr_selector3_4084;
wire[15:0] addr_remain3_4084;
address_decode_4 decoder_3_4084 = address_decode_4(addr_selector2_255[4],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4084,addr_remain3_4084);


wire[15:0] addr_selector3_4085;
wire[15:0] addr_remain3_4085;
address_decode_4 decoder_3_4085 = address_decode_4(addr_selector2_255[5],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4085,addr_remain3_4085);


wire[15:0] addr_selector3_4086;
wire[15:0] addr_remain3_4086;
address_decode_4 decoder_3_4086 = address_decode_4(addr_selector2_255[6],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4086,addr_remain3_4086);


wire[15:0] addr_selector3_4087;
wire[15:0] addr_remain3_4087;
address_decode_4 decoder_3_4087 = address_decode_4(addr_selector2_255[7],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4087,addr_remain3_4087);


wire[15:0] addr_selector3_4088;
wire[15:0] addr_remain3_4088;
address_decode_4 decoder_3_4088 = address_decode_4(addr_selector2_255[8],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4088,addr_remain3_4088);


wire[15:0] addr_selector3_4089;
wire[15:0] addr_remain3_4089;
address_decode_4 decoder_3_4089 = address_decode_4(addr_selector2_255[9],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4089,addr_remain3_4089);


wire[15:0] addr_selector3_4090;
wire[15:0] addr_remain3_4090;
address_decode_4 decoder_3_4090 = address_decode_4(addr_selector2_255[10],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4090,addr_remain3_4090);


wire[15:0] addr_selector3_4091;
wire[15:0] addr_remain3_4091;
address_decode_4 decoder_3_4091 = address_decode_4(addr_selector2_255[11],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4091,addr_remain3_4091);


wire[15:0] addr_selector3_4092;
wire[15:0] addr_remain3_4092;
address_decode_4 decoder_3_4092 = address_decode_4(addr_selector2_255[12],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4092,addr_remain3_4092);


wire[15:0] addr_selector3_4093;
wire[15:0] addr_remain3_4093;
address_decode_4 decoder_3_4093 = address_decode_4(addr_selector2_255[13],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4093,addr_remain3_4093);


wire[15:0] addr_selector3_4094;
wire[15:0] addr_remain3_4094;
address_decode_4 decoder_3_4094 = address_decode_4(addr_selector2_255[14],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4094,addr_remain3_4094);


wire[15:0] addr_selector3_4095;
wire[15:0] addr_remain3_4095;
address_decode_4 decoder_3_4095 = address_decode_4(addr_selector2_255[15],addr_remain2_255[15:0],addr_remain2_255,addr_selector3_4095,addr_remain3_4095);




assign addr_selector = {addr_selector3_0,addr_selector3_1,addr_selector3_2,addr_selector3_3,addr_selector3_4,addr_selector3_5,addr_selector3_6,addr_selector3_7,addr_selector3_8,addr_selector3_9,addr_selector3_10,addr_selector3_11,addr_selector3_12,addr_selector3_13,addr_selector3_14,addr_selector3_15,addr_selector3_16,addr_selector3_17,addr_selector3_18,addr_selector3_19,addr_selector3_20,addr_selector3_21,addr_selector3_22,addr_selector3_23,addr_selector3_24,addr_selector3_25,addr_selector3_26,addr_selector3_27,addr_selector3_28,addr_selector3_29,addr_selector3_30,addr_selector3_31,addr_selector3_32,addr_selector3_33,addr_selector3_34,addr_selector3_35,addr_selector3_36,addr_selector3_37,addr_selector3_38,addr_selector3_39,addr_selector3_40,addr_selector3_41,addr_selector3_42,addr_selector3_43,addr_selector3_44,addr_selector3_45,addr_selector3_46,addr_selector3_47,addr_selector3_48,addr_selector3_49,addr_selector3_50,addr_selector3_51,addr_selector3_52,addr_selector3_53,addr_selector3_54,addr_selector3_55,addr_selector3_56,addr_selector3_57,addr_selector3_58,addr_selector3_59,addr_selector3_60,addr_selector3_61,addr_selector3_62,addr_selector3_63,addr_selector3_64,addr_selector3_65,addr_selector3_66,addr_selector3_67,addr_selector3_68,addr_selector3_69,addr_selector3_70,addr_selector3_71,addr_selector3_72,addr_selector3_73,addr_selector3_74,addr_selector3_75,addr_selector3_76,addr_selector3_77,addr_selector3_78,addr_selector3_79,addr_selector3_80,addr_selector3_81,addr_selector3_82,addr_selector3_83,addr_selector3_84,addr_selector3_85,addr_selector3_86,addr_selector3_87,addr_selector3_88,addr_selector3_89,addr_selector3_90,addr_selector3_91,addr_selector3_92,addr_selector3_93,addr_selector3_94,addr_selector3_95,addr_selector3_96,addr_selector3_97,addr_selector3_98,addr_selector3_99,addr_selector3_100,addr_selector3_101,addr_selector3_102,addr_selector3_103,addr_selector3_104,addr_selector3_105,addr_selector3_106,addr_selector3_107,addr_selector3_108,addr_selector3_109,addr_selector3_110,addr_selector3_111,addr_selector3_112,addr_selector3_113,addr_selector3_114,addr_selector3_115,addr_selector3_116,addr_selector3_117,addr_selector3_118,addr_selector3_119,addr_selector3_120,addr_selector3_121,addr_selector3_122,addr_selector3_123,addr_selector3_124,addr_selector3_125,addr_selector3_126,addr_selector3_127,addr_selector3_128,addr_selector3_129,addr_selector3_130,addr_selector3_131,addr_selector3_132,addr_selector3_133,addr_selector3_134,addr_selector3_135,addr_selector3_136,addr_selector3_137,addr_selector3_138,addr_selector3_139,addr_selector3_140,addr_selector3_141,addr_selector3_142,addr_selector3_143,addr_selector3_144,addr_selector3_145,addr_selector3_146,addr_selector3_147,addr_selector3_148,addr_selector3_149,addr_selector3_150,addr_selector3_151,addr_selector3_152,addr_selector3_153,addr_selector3_154,addr_selector3_155,addr_selector3_156,addr_selector3_157,addr_selector3_158,addr_selector3_159,addr_selector3_160,addr_selector3_161,addr_selector3_162,addr_selector3_163,addr_selector3_164,addr_selector3_165,addr_selector3_166,addr_selector3_167,addr_selector3_168,addr_selector3_169,addr_selector3_170,addr_selector3_171,addr_selector3_172,addr_selector3_173,addr_selector3_174,addr_selector3_175,addr_selector3_176,addr_selector3_177,addr_selector3_178,addr_selector3_179,addr_selector3_180,addr_selector3_181,addr_selector3_182,addr_selector3_183,addr_selector3_184,addr_selector3_185,addr_selector3_186,addr_selector3_187,addr_selector3_188,addr_selector3_189,addr_selector3_190,addr_selector3_191,addr_selector3_192,addr_selector3_193,addr_selector3_194,addr_selector3_195,addr_selector3_196,addr_selector3_197,addr_selector3_198,addr_selector3_199,addr_selector3_200,addr_selector3_201,addr_selector3_202,addr_selector3_203,addr_selector3_204,addr_selector3_205,addr_selector3_206,addr_selector3_207,addr_selector3_208,addr_selector3_209,addr_selector3_210,addr_selector3_211,addr_selector3_212,addr_selector3_213,addr_selector3_214,addr_selector3_215,addr_selector3_216,addr_selector3_217,addr_selector3_218,addr_selector3_219,addr_selector3_220,addr_selector3_221,addr_selector3_222,addr_selector3_223,addr_selector3_224,addr_selector3_225,addr_selector3_226,addr_selector3_227,addr_selector3_228,addr_selector3_229,addr_selector3_230,addr_selector3_231,addr_selector3_232,addr_selector3_233,addr_selector3_234,addr_selector3_235,addr_selector3_236,addr_selector3_237,addr_selector3_238,addr_selector3_239,addr_selector3_240,addr_selector3_241,addr_selector3_242,addr_selector3_243,addr_selector3_244,addr_selector3_245,addr_selector3_246,addr_selector3_247,addr_selector3_248,addr_selector3_249,addr_selector3_250,addr_selector3_251,addr_selector3_252,addr_selector3_253,addr_selector3_254,addr_selector3_255,addr_selector3_256,addr_selector3_257,addr_selector3_258,addr_selector3_259,addr_selector3_260,addr_selector3_261,addr_selector3_262,addr_selector3_263,addr_selector3_264,addr_selector3_265,addr_selector3_266,addr_selector3_267,addr_selector3_268,addr_selector3_269,addr_selector3_270,addr_selector3_271,addr_selector3_272,addr_selector3_273,addr_selector3_274,addr_selector3_275,addr_selector3_276,addr_selector3_277,addr_selector3_278,addr_selector3_279,addr_selector3_280,addr_selector3_281,addr_selector3_282,addr_selector3_283,addr_selector3_284,addr_selector3_285,addr_selector3_286,addr_selector3_287,addr_selector3_288,addr_selector3_289,addr_selector3_290,addr_selector3_291,addr_selector3_292,addr_selector3_293,addr_selector3_294,addr_selector3_295,addr_selector3_296,addr_selector3_297,addr_selector3_298,addr_selector3_299,addr_selector3_300,addr_selector3_301,addr_selector3_302,addr_selector3_303,addr_selector3_304,addr_selector3_305,addr_selector3_306,addr_selector3_307,addr_selector3_308,addr_selector3_309,addr_selector3_310,addr_selector3_311,addr_selector3_312,addr_selector3_313,addr_selector3_314,addr_selector3_315,addr_selector3_316,addr_selector3_317,addr_selector3_318,addr_selector3_319,addr_selector3_320,addr_selector3_321,addr_selector3_322,addr_selector3_323,addr_selector3_324,addr_selector3_325,addr_selector3_326,addr_selector3_327,addr_selector3_328,addr_selector3_329,addr_selector3_330,addr_selector3_331,addr_selector3_332,addr_selector3_333,addr_selector3_334,addr_selector3_335,addr_selector3_336,addr_selector3_337,addr_selector3_338,addr_selector3_339,addr_selector3_340,addr_selector3_341,addr_selector3_342,addr_selector3_343,addr_selector3_344,addr_selector3_345,addr_selector3_346,addr_selector3_347,addr_selector3_348,addr_selector3_349,addr_selector3_350,addr_selector3_351,addr_selector3_352,addr_selector3_353,addr_selector3_354,addr_selector3_355,addr_selector3_356,addr_selector3_357,addr_selector3_358,addr_selector3_359,addr_selector3_360,addr_selector3_361,addr_selector3_362,addr_selector3_363,addr_selector3_364,addr_selector3_365,addr_selector3_366,addr_selector3_367,addr_selector3_368,addr_selector3_369,addr_selector3_370,addr_selector3_371,addr_selector3_372,addr_selector3_373,addr_selector3_374,addr_selector3_375,addr_selector3_376,addr_selector3_377,addr_selector3_378,addr_selector3_379,addr_selector3_380,addr_selector3_381,addr_selector3_382,addr_selector3_383,addr_selector3_384,addr_selector3_385,addr_selector3_386,addr_selector3_387,addr_selector3_388,addr_selector3_389,addr_selector3_390,addr_selector3_391,addr_selector3_392,addr_selector3_393,addr_selector3_394,addr_selector3_395,addr_selector3_396,addr_selector3_397,addr_selector3_398,addr_selector3_399,addr_selector3_400,addr_selector3_401,addr_selector3_402,addr_selector3_403,addr_selector3_404,addr_selector3_405,addr_selector3_406,addr_selector3_407,addr_selector3_408,addr_selector3_409,addr_selector3_410,addr_selector3_411,addr_selector3_412,addr_selector3_413,addr_selector3_414,addr_selector3_415,addr_selector3_416,addr_selector3_417,addr_selector3_418,addr_selector3_419,addr_selector3_420,addr_selector3_421,addr_selector3_422,addr_selector3_423,addr_selector3_424,addr_selector3_425,addr_selector3_426,addr_selector3_427,addr_selector3_428,addr_selector3_429,addr_selector3_430,addr_selector3_431,addr_selector3_432,addr_selector3_433,addr_selector3_434,addr_selector3_435,addr_selector3_436,addr_selector3_437,addr_selector3_438,addr_selector3_439,addr_selector3_440,addr_selector3_441,addr_selector3_442,addr_selector3_443,addr_selector3_444,addr_selector3_445,addr_selector3_446,addr_selector3_447,addr_selector3_448,addr_selector3_449,addr_selector3_450,addr_selector3_451,addr_selector3_452,addr_selector3_453,addr_selector3_454,addr_selector3_455,addr_selector3_456,addr_selector3_457,addr_selector3_458,addr_selector3_459,addr_selector3_460,addr_selector3_461,addr_selector3_462,addr_selector3_463,addr_selector3_464,addr_selector3_465,addr_selector3_466,addr_selector3_467,addr_selector3_468,addr_selector3_469,addr_selector3_470,addr_selector3_471,addr_selector3_472,addr_selector3_473,addr_selector3_474,addr_selector3_475,addr_selector3_476,addr_selector3_477,addr_selector3_478,addr_selector3_479,addr_selector3_480,addr_selector3_481,addr_selector3_482,addr_selector3_483,addr_selector3_484,addr_selector3_485,addr_selector3_486,addr_selector3_487,addr_selector3_488,addr_selector3_489,addr_selector3_490,addr_selector3_491,addr_selector3_492,addr_selector3_493,addr_selector3_494,addr_selector3_495,addr_selector3_496,addr_selector3_497,addr_selector3_498,addr_selector3_499,addr_selector3_500,addr_selector3_501,addr_selector3_502,addr_selector3_503,addr_selector3_504,addr_selector3_505,addr_selector3_506,addr_selector3_507,addr_selector3_508,addr_selector3_509,addr_selector3_510,addr_selector3_511,addr_selector3_512,addr_selector3_513,addr_selector3_514,addr_selector3_515,addr_selector3_516,addr_selector3_517,addr_selector3_518,addr_selector3_519,addr_selector3_520,addr_selector3_521,addr_selector3_522,addr_selector3_523,addr_selector3_524,addr_selector3_525,addr_selector3_526,addr_selector3_527,addr_selector3_528,addr_selector3_529,addr_selector3_530,addr_selector3_531,addr_selector3_532,addr_selector3_533,addr_selector3_534,addr_selector3_535,addr_selector3_536,addr_selector3_537,addr_selector3_538,addr_selector3_539,addr_selector3_540,addr_selector3_541,addr_selector3_542,addr_selector3_543,addr_selector3_544,addr_selector3_545,addr_selector3_546,addr_selector3_547,addr_selector3_548,addr_selector3_549,addr_selector3_550,addr_selector3_551,addr_selector3_552,addr_selector3_553,addr_selector3_554,addr_selector3_555,addr_selector3_556,addr_selector3_557,addr_selector3_558,addr_selector3_559,addr_selector3_560,addr_selector3_561,addr_selector3_562,addr_selector3_563,addr_selector3_564,addr_selector3_565,addr_selector3_566,addr_selector3_567,addr_selector3_568,addr_selector3_569,addr_selector3_570,addr_selector3_571,addr_selector3_572,addr_selector3_573,addr_selector3_574,addr_selector3_575,addr_selector3_576,addr_selector3_577,addr_selector3_578,addr_selector3_579,addr_selector3_580,addr_selector3_581,addr_selector3_582,addr_selector3_583,addr_selector3_584,addr_selector3_585,addr_selector3_586,addr_selector3_587,addr_selector3_588,addr_selector3_589,addr_selector3_590,addr_selector3_591,addr_selector3_592,addr_selector3_593,addr_selector3_594,addr_selector3_595,addr_selector3_596,addr_selector3_597,addr_selector3_598,addr_selector3_599,addr_selector3_600,addr_selector3_601,addr_selector3_602,addr_selector3_603,addr_selector3_604,addr_selector3_605,addr_selector3_606,addr_selector3_607,addr_selector3_608,addr_selector3_609,addr_selector3_610,addr_selector3_611,addr_selector3_612,addr_selector3_613,addr_selector3_614,addr_selector3_615,addr_selector3_616,addr_selector3_617,addr_selector3_618,addr_selector3_619,addr_selector3_620,addr_selector3_621,addr_selector3_622,addr_selector3_623,addr_selector3_624,addr_selector3_625,addr_selector3_626,addr_selector3_627,addr_selector3_628,addr_selector3_629,addr_selector3_630,addr_selector3_631,addr_selector3_632,addr_selector3_633,addr_selector3_634,addr_selector3_635,addr_selector3_636,addr_selector3_637,addr_selector3_638,addr_selector3_639,addr_selector3_640,addr_selector3_641,addr_selector3_642,addr_selector3_643,addr_selector3_644,addr_selector3_645,addr_selector3_646,addr_selector3_647,addr_selector3_648,addr_selector3_649,addr_selector3_650,addr_selector3_651,addr_selector3_652,addr_selector3_653,addr_selector3_654,addr_selector3_655,addr_selector3_656,addr_selector3_657,addr_selector3_658,addr_selector3_659,addr_selector3_660,addr_selector3_661,addr_selector3_662,addr_selector3_663,addr_selector3_664,addr_selector3_665,addr_selector3_666,addr_selector3_667,addr_selector3_668,addr_selector3_669,addr_selector3_670,addr_selector3_671,addr_selector3_672,addr_selector3_673,addr_selector3_674,addr_selector3_675,addr_selector3_676,addr_selector3_677,addr_selector3_678,addr_selector3_679,addr_selector3_680,addr_selector3_681,addr_selector3_682,addr_selector3_683,addr_selector3_684,addr_selector3_685,addr_selector3_686,addr_selector3_687,addr_selector3_688,addr_selector3_689,addr_selector3_690,addr_selector3_691,addr_selector3_692,addr_selector3_693,addr_selector3_694,addr_selector3_695,addr_selector3_696,addr_selector3_697,addr_selector3_698,addr_selector3_699,addr_selector3_700,addr_selector3_701,addr_selector3_702,addr_selector3_703,addr_selector3_704,addr_selector3_705,addr_selector3_706,addr_selector3_707,addr_selector3_708,addr_selector3_709,addr_selector3_710,addr_selector3_711,addr_selector3_712,addr_selector3_713,addr_selector3_714,addr_selector3_715,addr_selector3_716,addr_selector3_717,addr_selector3_718,addr_selector3_719,addr_selector3_720,addr_selector3_721,addr_selector3_722,addr_selector3_723,addr_selector3_724,addr_selector3_725,addr_selector3_726,addr_selector3_727,addr_selector3_728,addr_selector3_729,addr_selector3_730,addr_selector3_731,addr_selector3_732,addr_selector3_733,addr_selector3_734,addr_selector3_735,addr_selector3_736,addr_selector3_737,addr_selector3_738,addr_selector3_739,addr_selector3_740,addr_selector3_741,addr_selector3_742,addr_selector3_743,addr_selector3_744,addr_selector3_745,addr_selector3_746,addr_selector3_747,addr_selector3_748,addr_selector3_749,addr_selector3_750,addr_selector3_751,addr_selector3_752,addr_selector3_753,addr_selector3_754,addr_selector3_755,addr_selector3_756,addr_selector3_757,addr_selector3_758,addr_selector3_759,addr_selector3_760,addr_selector3_761,addr_selector3_762,addr_selector3_763,addr_selector3_764,addr_selector3_765,addr_selector3_766,addr_selector3_767,addr_selector3_768,addr_selector3_769,addr_selector3_770,addr_selector3_771,addr_selector3_772,addr_selector3_773,addr_selector3_774,addr_selector3_775,addr_selector3_776,addr_selector3_777,addr_selector3_778,addr_selector3_779,addr_selector3_780,addr_selector3_781,addr_selector3_782,addr_selector3_783,addr_selector3_784,addr_selector3_785,addr_selector3_786,addr_selector3_787,addr_selector3_788,addr_selector3_789,addr_selector3_790,addr_selector3_791,addr_selector3_792,addr_selector3_793,addr_selector3_794,addr_selector3_795,addr_selector3_796,addr_selector3_797,addr_selector3_798,addr_selector3_799,addr_selector3_800,addr_selector3_801,addr_selector3_802,addr_selector3_803,addr_selector3_804,addr_selector3_805,addr_selector3_806,addr_selector3_807,addr_selector3_808,addr_selector3_809,addr_selector3_810,addr_selector3_811,addr_selector3_812,addr_selector3_813,addr_selector3_814,addr_selector3_815,addr_selector3_816,addr_selector3_817,addr_selector3_818,addr_selector3_819,addr_selector3_820,addr_selector3_821,addr_selector3_822,addr_selector3_823,addr_selector3_824,addr_selector3_825,addr_selector3_826,addr_selector3_827,addr_selector3_828,addr_selector3_829,addr_selector3_830,addr_selector3_831,addr_selector3_832,addr_selector3_833,addr_selector3_834,addr_selector3_835,addr_selector3_836,addr_selector3_837,addr_selector3_838,addr_selector3_839,addr_selector3_840,addr_selector3_841,addr_selector3_842,addr_selector3_843,addr_selector3_844,addr_selector3_845,addr_selector3_846,addr_selector3_847,addr_selector3_848,addr_selector3_849,addr_selector3_850,addr_selector3_851,addr_selector3_852,addr_selector3_853,addr_selector3_854,addr_selector3_855,addr_selector3_856,addr_selector3_857,addr_selector3_858,addr_selector3_859,addr_selector3_860,addr_selector3_861,addr_selector3_862,addr_selector3_863,addr_selector3_864,addr_selector3_865,addr_selector3_866,addr_selector3_867,addr_selector3_868,addr_selector3_869,addr_selector3_870,addr_selector3_871,addr_selector3_872,addr_selector3_873,addr_selector3_874,addr_selector3_875,addr_selector3_876,addr_selector3_877,addr_selector3_878,addr_selector3_879,addr_selector3_880,addr_selector3_881,addr_selector3_882,addr_selector3_883,addr_selector3_884,addr_selector3_885,addr_selector3_886,addr_selector3_887,addr_selector3_888,addr_selector3_889,addr_selector3_890,addr_selector3_891,addr_selector3_892,addr_selector3_893,addr_selector3_894,addr_selector3_895,addr_selector3_896,addr_selector3_897,addr_selector3_898,addr_selector3_899,addr_selector3_900,addr_selector3_901,addr_selector3_902,addr_selector3_903,addr_selector3_904,addr_selector3_905,addr_selector3_906,addr_selector3_907,addr_selector3_908,addr_selector3_909,addr_selector3_910,addr_selector3_911,addr_selector3_912,addr_selector3_913,addr_selector3_914,addr_selector3_915,addr_selector3_916,addr_selector3_917,addr_selector3_918,addr_selector3_919,addr_selector3_920,addr_selector3_921,addr_selector3_922,addr_selector3_923,addr_selector3_924,addr_selector3_925,addr_selector3_926,addr_selector3_927,addr_selector3_928,addr_selector3_929,addr_selector3_930,addr_selector3_931,addr_selector3_932,addr_selector3_933,addr_selector3_934,addr_selector3_935,addr_selector3_936,addr_selector3_937,addr_selector3_938,addr_selector3_939,addr_selector3_940,addr_selector3_941,addr_selector3_942,addr_selector3_943,addr_selector3_944,addr_selector3_945,addr_selector3_946,addr_selector3_947,addr_selector3_948,addr_selector3_949,addr_selector3_950,addr_selector3_951,addr_selector3_952,addr_selector3_953,addr_selector3_954,addr_selector3_955,addr_selector3_956,addr_selector3_957,addr_selector3_958,addr_selector3_959,addr_selector3_960,addr_selector3_961,addr_selector3_962,addr_selector3_963,addr_selector3_964,addr_selector3_965,addr_selector3_966,addr_selector3_967,addr_selector3_968,addr_selector3_969,addr_selector3_970,addr_selector3_971,addr_selector3_972,addr_selector3_973,addr_selector3_974,addr_selector3_975,addr_selector3_976,addr_selector3_977,addr_selector3_978,addr_selector3_979,addr_selector3_980,addr_selector3_981,addr_selector3_982,addr_selector3_983,addr_selector3_984,addr_selector3_985,addr_selector3_986,addr_selector3_987,addr_selector3_988,addr_selector3_989,addr_selector3_990,addr_selector3_991,addr_selector3_992,addr_selector3_993,addr_selector3_994,addr_selector3_995,addr_selector3_996,addr_selector3_997,addr_selector3_998,addr_selector3_999,addr_selector3_1000,addr_selector3_1001,addr_selector3_1002,addr_selector3_1003,addr_selector3_1004,addr_selector3_1005,addr_selector3_1006,addr_selector3_1007,addr_selector3_1008,addr_selector3_1009,addr_selector3_1010,addr_selector3_1011,addr_selector3_1012,addr_selector3_1013,addr_selector3_1014,addr_selector3_1015,addr_selector3_1016,addr_selector3_1017,addr_selector3_1018,addr_selector3_1019,addr_selector3_1020,addr_selector3_1021,addr_selector3_1022,addr_selector3_1023,addr_selector3_1024,addr_selector3_1025,addr_selector3_1026,addr_selector3_1027,addr_selector3_1028,addr_selector3_1029,addr_selector3_1030,addr_selector3_1031,addr_selector3_1032,addr_selector3_1033,addr_selector3_1034,addr_selector3_1035,addr_selector3_1036,addr_selector3_1037,addr_selector3_1038,addr_selector3_1039,addr_selector3_1040,addr_selector3_1041,addr_selector3_1042,addr_selector3_1043,addr_selector3_1044,addr_selector3_1045,addr_selector3_1046,addr_selector3_1047,addr_selector3_1048,addr_selector3_1049,addr_selector3_1050,addr_selector3_1051,addr_selector3_1052,addr_selector3_1053,addr_selector3_1054,addr_selector3_1055,addr_selector3_1056,addr_selector3_1057,addr_selector3_1058,addr_selector3_1059,addr_selector3_1060,addr_selector3_1061,addr_selector3_1062,addr_selector3_1063,addr_selector3_1064,addr_selector3_1065,addr_selector3_1066,addr_selector3_1067,addr_selector3_1068,addr_selector3_1069,addr_selector3_1070,addr_selector3_1071,addr_selector3_1072,addr_selector3_1073,addr_selector3_1074,addr_selector3_1075,addr_selector3_1076,addr_selector3_1077,addr_selector3_1078,addr_selector3_1079,addr_selector3_1080,addr_selector3_1081,addr_selector3_1082,addr_selector3_1083,addr_selector3_1084,addr_selector3_1085,addr_selector3_1086,addr_selector3_1087,addr_selector3_1088,addr_selector3_1089,addr_selector3_1090,addr_selector3_1091,addr_selector3_1092,addr_selector3_1093,addr_selector3_1094,addr_selector3_1095,addr_selector3_1096,addr_selector3_1097,addr_selector3_1098,addr_selector3_1099,addr_selector3_1100,addr_selector3_1101,addr_selector3_1102,addr_selector3_1103,addr_selector3_1104,addr_selector3_1105,addr_selector3_1106,addr_selector3_1107,addr_selector3_1108,addr_selector3_1109,addr_selector3_1110,addr_selector3_1111,addr_selector3_1112,addr_selector3_1113,addr_selector3_1114,addr_selector3_1115,addr_selector3_1116,addr_selector3_1117,addr_selector3_1118,addr_selector3_1119,addr_selector3_1120,addr_selector3_1121,addr_selector3_1122,addr_selector3_1123,addr_selector3_1124,addr_selector3_1125,addr_selector3_1126,addr_selector3_1127,addr_selector3_1128,addr_selector3_1129,addr_selector3_1130,addr_selector3_1131,addr_selector3_1132,addr_selector3_1133,addr_selector3_1134,addr_selector3_1135,addr_selector3_1136,addr_selector3_1137,addr_selector3_1138,addr_selector3_1139,addr_selector3_1140,addr_selector3_1141,addr_selector3_1142,addr_selector3_1143,addr_selector3_1144,addr_selector3_1145,addr_selector3_1146,addr_selector3_1147,addr_selector3_1148,addr_selector3_1149,addr_selector3_1150,addr_selector3_1151,addr_selector3_1152,addr_selector3_1153,addr_selector3_1154,addr_selector3_1155,addr_selector3_1156,addr_selector3_1157,addr_selector3_1158,addr_selector3_1159,addr_selector3_1160,addr_selector3_1161,addr_selector3_1162,addr_selector3_1163,addr_selector3_1164,addr_selector3_1165,addr_selector3_1166,addr_selector3_1167,addr_selector3_1168,addr_selector3_1169,addr_selector3_1170,addr_selector3_1171,addr_selector3_1172,addr_selector3_1173,addr_selector3_1174,addr_selector3_1175,addr_selector3_1176,addr_selector3_1177,addr_selector3_1178,addr_selector3_1179,addr_selector3_1180,addr_selector3_1181,addr_selector3_1182,addr_selector3_1183,addr_selector3_1184,addr_selector3_1185,addr_selector3_1186,addr_selector3_1187,addr_selector3_1188,addr_selector3_1189,addr_selector3_1190,addr_selector3_1191,addr_selector3_1192,addr_selector3_1193,addr_selector3_1194,addr_selector3_1195,addr_selector3_1196,addr_selector3_1197,addr_selector3_1198,addr_selector3_1199,addr_selector3_1200,addr_selector3_1201,addr_selector3_1202,addr_selector3_1203,addr_selector3_1204,addr_selector3_1205,addr_selector3_1206,addr_selector3_1207,addr_selector3_1208,addr_selector3_1209,addr_selector3_1210,addr_selector3_1211,addr_selector3_1212,addr_selector3_1213,addr_selector3_1214,addr_selector3_1215,addr_selector3_1216,addr_selector3_1217,addr_selector3_1218,addr_selector3_1219,addr_selector3_1220,addr_selector3_1221,addr_selector3_1222,addr_selector3_1223,addr_selector3_1224,addr_selector3_1225,addr_selector3_1226,addr_selector3_1227,addr_selector3_1228,addr_selector3_1229,addr_selector3_1230,addr_selector3_1231,addr_selector3_1232,addr_selector3_1233,addr_selector3_1234,addr_selector3_1235,addr_selector3_1236,addr_selector3_1237,addr_selector3_1238,addr_selector3_1239,addr_selector3_1240,addr_selector3_1241,addr_selector3_1242,addr_selector3_1243,addr_selector3_1244,addr_selector3_1245,addr_selector3_1246,addr_selector3_1247,addr_selector3_1248,addr_selector3_1249,addr_selector3_1250,addr_selector3_1251,addr_selector3_1252,addr_selector3_1253,addr_selector3_1254,addr_selector3_1255,addr_selector3_1256,addr_selector3_1257,addr_selector3_1258,addr_selector3_1259,addr_selector3_1260,addr_selector3_1261,addr_selector3_1262,addr_selector3_1263,addr_selector3_1264,addr_selector3_1265,addr_selector3_1266,addr_selector3_1267,addr_selector3_1268,addr_selector3_1269,addr_selector3_1270,addr_selector3_1271,addr_selector3_1272,addr_selector3_1273,addr_selector3_1274,addr_selector3_1275,addr_selector3_1276,addr_selector3_1277,addr_selector3_1278,addr_selector3_1279,addr_selector3_1280,addr_selector3_1281,addr_selector3_1282,addr_selector3_1283,addr_selector3_1284,addr_selector3_1285,addr_selector3_1286,addr_selector3_1287,addr_selector3_1288,addr_selector3_1289,addr_selector3_1290,addr_selector3_1291,addr_selector3_1292,addr_selector3_1293,addr_selector3_1294,addr_selector3_1295,addr_selector3_1296,addr_selector3_1297,addr_selector3_1298,addr_selector3_1299,addr_selector3_1300,addr_selector3_1301,addr_selector3_1302,addr_selector3_1303,addr_selector3_1304,addr_selector3_1305,addr_selector3_1306,addr_selector3_1307,addr_selector3_1308,addr_selector3_1309,addr_selector3_1310,addr_selector3_1311,addr_selector3_1312,addr_selector3_1313,addr_selector3_1314,addr_selector3_1315,addr_selector3_1316,addr_selector3_1317,addr_selector3_1318,addr_selector3_1319,addr_selector3_1320,addr_selector3_1321,addr_selector3_1322,addr_selector3_1323,addr_selector3_1324,addr_selector3_1325,addr_selector3_1326,addr_selector3_1327,addr_selector3_1328,addr_selector3_1329,addr_selector3_1330,addr_selector3_1331,addr_selector3_1332,addr_selector3_1333,addr_selector3_1334,addr_selector3_1335,addr_selector3_1336,addr_selector3_1337,addr_selector3_1338,addr_selector3_1339,addr_selector3_1340,addr_selector3_1341,addr_selector3_1342,addr_selector3_1343,addr_selector3_1344,addr_selector3_1345,addr_selector3_1346,addr_selector3_1347,addr_selector3_1348,addr_selector3_1349,addr_selector3_1350,addr_selector3_1351,addr_selector3_1352,addr_selector3_1353,addr_selector3_1354,addr_selector3_1355,addr_selector3_1356,addr_selector3_1357,addr_selector3_1358,addr_selector3_1359,addr_selector3_1360,addr_selector3_1361,addr_selector3_1362,addr_selector3_1363,addr_selector3_1364,addr_selector3_1365,addr_selector3_1366,addr_selector3_1367,addr_selector3_1368,addr_selector3_1369,addr_selector3_1370,addr_selector3_1371,addr_selector3_1372,addr_selector3_1373,addr_selector3_1374,addr_selector3_1375,addr_selector3_1376,addr_selector3_1377,addr_selector3_1378,addr_selector3_1379,addr_selector3_1380,addr_selector3_1381,addr_selector3_1382,addr_selector3_1383,addr_selector3_1384,addr_selector3_1385,addr_selector3_1386,addr_selector3_1387,addr_selector3_1388,addr_selector3_1389,addr_selector3_1390,addr_selector3_1391,addr_selector3_1392,addr_selector3_1393,addr_selector3_1394,addr_selector3_1395,addr_selector3_1396,addr_selector3_1397,addr_selector3_1398,addr_selector3_1399,addr_selector3_1400,addr_selector3_1401,addr_selector3_1402,addr_selector3_1403,addr_selector3_1404,addr_selector3_1405,addr_selector3_1406,addr_selector3_1407,addr_selector3_1408,addr_selector3_1409,addr_selector3_1410,addr_selector3_1411,addr_selector3_1412,addr_selector3_1413,addr_selector3_1414,addr_selector3_1415,addr_selector3_1416,addr_selector3_1417,addr_selector3_1418,addr_selector3_1419,addr_selector3_1420,addr_selector3_1421,addr_selector3_1422,addr_selector3_1423,addr_selector3_1424,addr_selector3_1425,addr_selector3_1426,addr_selector3_1427,addr_selector3_1428,addr_selector3_1429,addr_selector3_1430,addr_selector3_1431,addr_selector3_1432,addr_selector3_1433,addr_selector3_1434,addr_selector3_1435,addr_selector3_1436,addr_selector3_1437,addr_selector3_1438,addr_selector3_1439,addr_selector3_1440,addr_selector3_1441,addr_selector3_1442,addr_selector3_1443,addr_selector3_1444,addr_selector3_1445,addr_selector3_1446,addr_selector3_1447,addr_selector3_1448,addr_selector3_1449,addr_selector3_1450,addr_selector3_1451,addr_selector3_1452,addr_selector3_1453,addr_selector3_1454,addr_selector3_1455,addr_selector3_1456,addr_selector3_1457,addr_selector3_1458,addr_selector3_1459,addr_selector3_1460,addr_selector3_1461,addr_selector3_1462,addr_selector3_1463,addr_selector3_1464,addr_selector3_1465,addr_selector3_1466,addr_selector3_1467,addr_selector3_1468,addr_selector3_1469,addr_selector3_1470,addr_selector3_1471,addr_selector3_1472,addr_selector3_1473,addr_selector3_1474,addr_selector3_1475,addr_selector3_1476,addr_selector3_1477,addr_selector3_1478,addr_selector3_1479,addr_selector3_1480,addr_selector3_1481,addr_selector3_1482,addr_selector3_1483,addr_selector3_1484,addr_selector3_1485,addr_selector3_1486,addr_selector3_1487,addr_selector3_1488,addr_selector3_1489,addr_selector3_1490,addr_selector3_1491,addr_selector3_1492,addr_selector3_1493,addr_selector3_1494,addr_selector3_1495,addr_selector3_1496,addr_selector3_1497,addr_selector3_1498,addr_selector3_1499,addr_selector3_1500,addr_selector3_1501,addr_selector3_1502,addr_selector3_1503,addr_selector3_1504,addr_selector3_1505,addr_selector3_1506,addr_selector3_1507,addr_selector3_1508,addr_selector3_1509,addr_selector3_1510,addr_selector3_1511,addr_selector3_1512,addr_selector3_1513,addr_selector3_1514,addr_selector3_1515,addr_selector3_1516,addr_selector3_1517,addr_selector3_1518,addr_selector3_1519,addr_selector3_1520,addr_selector3_1521,addr_selector3_1522,addr_selector3_1523,addr_selector3_1524,addr_selector3_1525,addr_selector3_1526,addr_selector3_1527,addr_selector3_1528,addr_selector3_1529,addr_selector3_1530,addr_selector3_1531,addr_selector3_1532,addr_selector3_1533,addr_selector3_1534,addr_selector3_1535,addr_selector3_1536,addr_selector3_1537,addr_selector3_1538,addr_selector3_1539,addr_selector3_1540,addr_selector3_1541,addr_selector3_1542,addr_selector3_1543,addr_selector3_1544,addr_selector3_1545,addr_selector3_1546,addr_selector3_1547,addr_selector3_1548,addr_selector3_1549,addr_selector3_1550,addr_selector3_1551,addr_selector3_1552,addr_selector3_1553,addr_selector3_1554,addr_selector3_1555,addr_selector3_1556,addr_selector3_1557,addr_selector3_1558,addr_selector3_1559,addr_selector3_1560,addr_selector3_1561,addr_selector3_1562,addr_selector3_1563,addr_selector3_1564,addr_selector3_1565,addr_selector3_1566,addr_selector3_1567,addr_selector3_1568,addr_selector3_1569,addr_selector3_1570,addr_selector3_1571,addr_selector3_1572,addr_selector3_1573,addr_selector3_1574,addr_selector3_1575,addr_selector3_1576,addr_selector3_1577,addr_selector3_1578,addr_selector3_1579,addr_selector3_1580,addr_selector3_1581,addr_selector3_1582,addr_selector3_1583,addr_selector3_1584,addr_selector3_1585,addr_selector3_1586,addr_selector3_1587,addr_selector3_1588,addr_selector3_1589,addr_selector3_1590,addr_selector3_1591,addr_selector3_1592,addr_selector3_1593,addr_selector3_1594,addr_selector3_1595,addr_selector3_1596,addr_selector3_1597,addr_selector3_1598,addr_selector3_1599,addr_selector3_1600,addr_selector3_1601,addr_selector3_1602,addr_selector3_1603,addr_selector3_1604,addr_selector3_1605,addr_selector3_1606,addr_selector3_1607,addr_selector3_1608,addr_selector3_1609,addr_selector3_1610,addr_selector3_1611,addr_selector3_1612,addr_selector3_1613,addr_selector3_1614,addr_selector3_1615,addr_selector3_1616,addr_selector3_1617,addr_selector3_1618,addr_selector3_1619,addr_selector3_1620,addr_selector3_1621,addr_selector3_1622,addr_selector3_1623,addr_selector3_1624,addr_selector3_1625,addr_selector3_1626,addr_selector3_1627,addr_selector3_1628,addr_selector3_1629,addr_selector3_1630,addr_selector3_1631,addr_selector3_1632,addr_selector3_1633,addr_selector3_1634,addr_selector3_1635,addr_selector3_1636,addr_selector3_1637,addr_selector3_1638,addr_selector3_1639,addr_selector3_1640,addr_selector3_1641,addr_selector3_1642,addr_selector3_1643,addr_selector3_1644,addr_selector3_1645,addr_selector3_1646,addr_selector3_1647,addr_selector3_1648,addr_selector3_1649,addr_selector3_1650,addr_selector3_1651,addr_selector3_1652,addr_selector3_1653,addr_selector3_1654,addr_selector3_1655,addr_selector3_1656,addr_selector3_1657,addr_selector3_1658,addr_selector3_1659,addr_selector3_1660,addr_selector3_1661,addr_selector3_1662,addr_selector3_1663,addr_selector3_1664,addr_selector3_1665,addr_selector3_1666,addr_selector3_1667,addr_selector3_1668,addr_selector3_1669,addr_selector3_1670,addr_selector3_1671,addr_selector3_1672,addr_selector3_1673,addr_selector3_1674,addr_selector3_1675,addr_selector3_1676,addr_selector3_1677,addr_selector3_1678,addr_selector3_1679,addr_selector3_1680,addr_selector3_1681,addr_selector3_1682,addr_selector3_1683,addr_selector3_1684,addr_selector3_1685,addr_selector3_1686,addr_selector3_1687,addr_selector3_1688,addr_selector3_1689,addr_selector3_1690,addr_selector3_1691,addr_selector3_1692,addr_selector3_1693,addr_selector3_1694,addr_selector3_1695,addr_selector3_1696,addr_selector3_1697,addr_selector3_1698,addr_selector3_1699,addr_selector3_1700,addr_selector3_1701,addr_selector3_1702,addr_selector3_1703,addr_selector3_1704,addr_selector3_1705,addr_selector3_1706,addr_selector3_1707,addr_selector3_1708,addr_selector3_1709,addr_selector3_1710,addr_selector3_1711,addr_selector3_1712,addr_selector3_1713,addr_selector3_1714,addr_selector3_1715,addr_selector3_1716,addr_selector3_1717,addr_selector3_1718,addr_selector3_1719,addr_selector3_1720,addr_selector3_1721,addr_selector3_1722,addr_selector3_1723,addr_selector3_1724,addr_selector3_1725,addr_selector3_1726,addr_selector3_1727,addr_selector3_1728,addr_selector3_1729,addr_selector3_1730,addr_selector3_1731,addr_selector3_1732,addr_selector3_1733,addr_selector3_1734,addr_selector3_1735,addr_selector3_1736,addr_selector3_1737,addr_selector3_1738,addr_selector3_1739,addr_selector3_1740,addr_selector3_1741,addr_selector3_1742,addr_selector3_1743,addr_selector3_1744,addr_selector3_1745,addr_selector3_1746,addr_selector3_1747,addr_selector3_1748,addr_selector3_1749,addr_selector3_1750,addr_selector3_1751,addr_selector3_1752,addr_selector3_1753,addr_selector3_1754,addr_selector3_1755,addr_selector3_1756,addr_selector3_1757,addr_selector3_1758,addr_selector3_1759,addr_selector3_1760,addr_selector3_1761,addr_selector3_1762,addr_selector3_1763,addr_selector3_1764,addr_selector3_1765,addr_selector3_1766,addr_selector3_1767,addr_selector3_1768,addr_selector3_1769,addr_selector3_1770,addr_selector3_1771,addr_selector3_1772,addr_selector3_1773,addr_selector3_1774,addr_selector3_1775,addr_selector3_1776,addr_selector3_1777,addr_selector3_1778,addr_selector3_1779,addr_selector3_1780,addr_selector3_1781,addr_selector3_1782,addr_selector3_1783,addr_selector3_1784,addr_selector3_1785,addr_selector3_1786,addr_selector3_1787,addr_selector3_1788,addr_selector3_1789,addr_selector3_1790,addr_selector3_1791,addr_selector3_1792,addr_selector3_1793,addr_selector3_1794,addr_selector3_1795,addr_selector3_1796,addr_selector3_1797,addr_selector3_1798,addr_selector3_1799,addr_selector3_1800,addr_selector3_1801,addr_selector3_1802,addr_selector3_1803,addr_selector3_1804,addr_selector3_1805,addr_selector3_1806,addr_selector3_1807,addr_selector3_1808,addr_selector3_1809,addr_selector3_1810,addr_selector3_1811,addr_selector3_1812,addr_selector3_1813,addr_selector3_1814,addr_selector3_1815,addr_selector3_1816,addr_selector3_1817,addr_selector3_1818,addr_selector3_1819,addr_selector3_1820,addr_selector3_1821,addr_selector3_1822,addr_selector3_1823,addr_selector3_1824,addr_selector3_1825,addr_selector3_1826,addr_selector3_1827,addr_selector3_1828,addr_selector3_1829,addr_selector3_1830,addr_selector3_1831,addr_selector3_1832,addr_selector3_1833,addr_selector3_1834,addr_selector3_1835,addr_selector3_1836,addr_selector3_1837,addr_selector3_1838,addr_selector3_1839,addr_selector3_1840,addr_selector3_1841,addr_selector3_1842,addr_selector3_1843,addr_selector3_1844,addr_selector3_1845,addr_selector3_1846,addr_selector3_1847,addr_selector3_1848,addr_selector3_1849,addr_selector3_1850,addr_selector3_1851,addr_selector3_1852,addr_selector3_1853,addr_selector3_1854,addr_selector3_1855,addr_selector3_1856,addr_selector3_1857,addr_selector3_1858,addr_selector3_1859,addr_selector3_1860,addr_selector3_1861,addr_selector3_1862,addr_selector3_1863,addr_selector3_1864,addr_selector3_1865,addr_selector3_1866,addr_selector3_1867,addr_selector3_1868,addr_selector3_1869,addr_selector3_1870,addr_selector3_1871,addr_selector3_1872,addr_selector3_1873,addr_selector3_1874,addr_selector3_1875,addr_selector3_1876,addr_selector3_1877,addr_selector3_1878,addr_selector3_1879,addr_selector3_1880,addr_selector3_1881,addr_selector3_1882,addr_selector3_1883,addr_selector3_1884,addr_selector3_1885,addr_selector3_1886,addr_selector3_1887,addr_selector3_1888,addr_selector3_1889,addr_selector3_1890,addr_selector3_1891,addr_selector3_1892,addr_selector3_1893,addr_selector3_1894,addr_selector3_1895,addr_selector3_1896,addr_selector3_1897,addr_selector3_1898,addr_selector3_1899,addr_selector3_1900,addr_selector3_1901,addr_selector3_1902,addr_selector3_1903,addr_selector3_1904,addr_selector3_1905,addr_selector3_1906,addr_selector3_1907,addr_selector3_1908,addr_selector3_1909,addr_selector3_1910,addr_selector3_1911,addr_selector3_1912,addr_selector3_1913,addr_selector3_1914,addr_selector3_1915,addr_selector3_1916,addr_selector3_1917,addr_selector3_1918,addr_selector3_1919,addr_selector3_1920,addr_selector3_1921,addr_selector3_1922,addr_selector3_1923,addr_selector3_1924,addr_selector3_1925,addr_selector3_1926,addr_selector3_1927,addr_selector3_1928,addr_selector3_1929,addr_selector3_1930,addr_selector3_1931,addr_selector3_1932,addr_selector3_1933,addr_selector3_1934,addr_selector3_1935,addr_selector3_1936,addr_selector3_1937,addr_selector3_1938,addr_selector3_1939,addr_selector3_1940,addr_selector3_1941,addr_selector3_1942,addr_selector3_1943,addr_selector3_1944,addr_selector3_1945,addr_selector3_1946,addr_selector3_1947,addr_selector3_1948,addr_selector3_1949,addr_selector3_1950,addr_selector3_1951,addr_selector3_1952,addr_selector3_1953,addr_selector3_1954,addr_selector3_1955,addr_selector3_1956,addr_selector3_1957,addr_selector3_1958,addr_selector3_1959,addr_selector3_1960,addr_selector3_1961,addr_selector3_1962,addr_selector3_1963,addr_selector3_1964,addr_selector3_1965,addr_selector3_1966,addr_selector3_1967,addr_selector3_1968,addr_selector3_1969,addr_selector3_1970,addr_selector3_1971,addr_selector3_1972,addr_selector3_1973,addr_selector3_1974,addr_selector3_1975,addr_selector3_1976,addr_selector3_1977,addr_selector3_1978,addr_selector3_1979,addr_selector3_1980,addr_selector3_1981,addr_selector3_1982,addr_selector3_1983,addr_selector3_1984,addr_selector3_1985,addr_selector3_1986,addr_selector3_1987,addr_selector3_1988,addr_selector3_1989,addr_selector3_1990,addr_selector3_1991,addr_selector3_1992,addr_selector3_1993,addr_selector3_1994,addr_selector3_1995,addr_selector3_1996,addr_selector3_1997,addr_selector3_1998,addr_selector3_1999,addr_selector3_2000,addr_selector3_2001,addr_selector3_2002,addr_selector3_2003,addr_selector3_2004,addr_selector3_2005,addr_selector3_2006,addr_selector3_2007,addr_selector3_2008,addr_selector3_2009,addr_selector3_2010,addr_selector3_2011,addr_selector3_2012,addr_selector3_2013,addr_selector3_2014,addr_selector3_2015,addr_selector3_2016,addr_selector3_2017,addr_selector3_2018,addr_selector3_2019,addr_selector3_2020,addr_selector3_2021,addr_selector3_2022,addr_selector3_2023,addr_selector3_2024,addr_selector3_2025,addr_selector3_2026,addr_selector3_2027,addr_selector3_2028,addr_selector3_2029,addr_selector3_2030,addr_selector3_2031,addr_selector3_2032,addr_selector3_2033,addr_selector3_2034,addr_selector3_2035,addr_selector3_2036,addr_selector3_2037,addr_selector3_2038,addr_selector3_2039,addr_selector3_2040,addr_selector3_2041,addr_selector3_2042,addr_selector3_2043,addr_selector3_2044,addr_selector3_2045,addr_selector3_2046,addr_selector3_2047,addr_selector3_2048,addr_selector3_2049,addr_selector3_2050,addr_selector3_2051,addr_selector3_2052,addr_selector3_2053,addr_selector3_2054,addr_selector3_2055,addr_selector3_2056,addr_selector3_2057,addr_selector3_2058,addr_selector3_2059,addr_selector3_2060,addr_selector3_2061,addr_selector3_2062,addr_selector3_2063,addr_selector3_2064,addr_selector3_2065,addr_selector3_2066,addr_selector3_2067,addr_selector3_2068,addr_selector3_2069,addr_selector3_2070,addr_selector3_2071,addr_selector3_2072,addr_selector3_2073,addr_selector3_2074,addr_selector3_2075,addr_selector3_2076,addr_selector3_2077,addr_selector3_2078,addr_selector3_2079,addr_selector3_2080,addr_selector3_2081,addr_selector3_2082,addr_selector3_2083,addr_selector3_2084,addr_selector3_2085,addr_selector3_2086,addr_selector3_2087,addr_selector3_2088,addr_selector3_2089,addr_selector3_2090,addr_selector3_2091,addr_selector3_2092,addr_selector3_2093,addr_selector3_2094,addr_selector3_2095,addr_selector3_2096,addr_selector3_2097,addr_selector3_2098,addr_selector3_2099,addr_selector3_2100,addr_selector3_2101,addr_selector3_2102,addr_selector3_2103,addr_selector3_2104,addr_selector3_2105,addr_selector3_2106,addr_selector3_2107,addr_selector3_2108,addr_selector3_2109,addr_selector3_2110,addr_selector3_2111,addr_selector3_2112,addr_selector3_2113,addr_selector3_2114,addr_selector3_2115,addr_selector3_2116,addr_selector3_2117,addr_selector3_2118,addr_selector3_2119,addr_selector3_2120,addr_selector3_2121,addr_selector3_2122,addr_selector3_2123,addr_selector3_2124,addr_selector3_2125,addr_selector3_2126,addr_selector3_2127,addr_selector3_2128,addr_selector3_2129,addr_selector3_2130,addr_selector3_2131,addr_selector3_2132,addr_selector3_2133,addr_selector3_2134,addr_selector3_2135,addr_selector3_2136,addr_selector3_2137,addr_selector3_2138,addr_selector3_2139,addr_selector3_2140,addr_selector3_2141,addr_selector3_2142,addr_selector3_2143,addr_selector3_2144,addr_selector3_2145,addr_selector3_2146,addr_selector3_2147,addr_selector3_2148,addr_selector3_2149,addr_selector3_2150,addr_selector3_2151,addr_selector3_2152,addr_selector3_2153,addr_selector3_2154,addr_selector3_2155,addr_selector3_2156,addr_selector3_2157,addr_selector3_2158,addr_selector3_2159,addr_selector3_2160,addr_selector3_2161,addr_selector3_2162,addr_selector3_2163,addr_selector3_2164,addr_selector3_2165,addr_selector3_2166,addr_selector3_2167,addr_selector3_2168,addr_selector3_2169,addr_selector3_2170,addr_selector3_2171,addr_selector3_2172,addr_selector3_2173,addr_selector3_2174,addr_selector3_2175,addr_selector3_2176,addr_selector3_2177,addr_selector3_2178,addr_selector3_2179,addr_selector3_2180,addr_selector3_2181,addr_selector3_2182,addr_selector3_2183,addr_selector3_2184,addr_selector3_2185,addr_selector3_2186,addr_selector3_2187,addr_selector3_2188,addr_selector3_2189,addr_selector3_2190,addr_selector3_2191,addr_selector3_2192,addr_selector3_2193,addr_selector3_2194,addr_selector3_2195,addr_selector3_2196,addr_selector3_2197,addr_selector3_2198,addr_selector3_2199,addr_selector3_2200,addr_selector3_2201,addr_selector3_2202,addr_selector3_2203,addr_selector3_2204,addr_selector3_2205,addr_selector3_2206,addr_selector3_2207,addr_selector3_2208,addr_selector3_2209,addr_selector3_2210,addr_selector3_2211,addr_selector3_2212,addr_selector3_2213,addr_selector3_2214,addr_selector3_2215,addr_selector3_2216,addr_selector3_2217,addr_selector3_2218,addr_selector3_2219,addr_selector3_2220,addr_selector3_2221,addr_selector3_2222,addr_selector3_2223,addr_selector3_2224,addr_selector3_2225,addr_selector3_2226,addr_selector3_2227,addr_selector3_2228,addr_selector3_2229,addr_selector3_2230,addr_selector3_2231,addr_selector3_2232,addr_selector3_2233,addr_selector3_2234,addr_selector3_2235,addr_selector3_2236,addr_selector3_2237,addr_selector3_2238,addr_selector3_2239,addr_selector3_2240,addr_selector3_2241,addr_selector3_2242,addr_selector3_2243,addr_selector3_2244,addr_selector3_2245,addr_selector3_2246,addr_selector3_2247,addr_selector3_2248,addr_selector3_2249,addr_selector3_2250,addr_selector3_2251,addr_selector3_2252,addr_selector3_2253,addr_selector3_2254,addr_selector3_2255,addr_selector3_2256,addr_selector3_2257,addr_selector3_2258,addr_selector3_2259,addr_selector3_2260,addr_selector3_2261,addr_selector3_2262,addr_selector3_2263,addr_selector3_2264,addr_selector3_2265,addr_selector3_2266,addr_selector3_2267,addr_selector3_2268,addr_selector3_2269,addr_selector3_2270,addr_selector3_2271,addr_selector3_2272,addr_selector3_2273,addr_selector3_2274,addr_selector3_2275,addr_selector3_2276,addr_selector3_2277,addr_selector3_2278,addr_selector3_2279,addr_selector3_2280,addr_selector3_2281,addr_selector3_2282,addr_selector3_2283,addr_selector3_2284,addr_selector3_2285,addr_selector3_2286,addr_selector3_2287,addr_selector3_2288,addr_selector3_2289,addr_selector3_2290,addr_selector3_2291,addr_selector3_2292,addr_selector3_2293,addr_selector3_2294,addr_selector3_2295,addr_selector3_2296,addr_selector3_2297,addr_selector3_2298,addr_selector3_2299,addr_selector3_2300,addr_selector3_2301,addr_selector3_2302,addr_selector3_2303,addr_selector3_2304,addr_selector3_2305,addr_selector3_2306,addr_selector3_2307,addr_selector3_2308,addr_selector3_2309,addr_selector3_2310,addr_selector3_2311,addr_selector3_2312,addr_selector3_2313,addr_selector3_2314,addr_selector3_2315,addr_selector3_2316,addr_selector3_2317,addr_selector3_2318,addr_selector3_2319,addr_selector3_2320,addr_selector3_2321,addr_selector3_2322,addr_selector3_2323,addr_selector3_2324,addr_selector3_2325,addr_selector3_2326,addr_selector3_2327,addr_selector3_2328,addr_selector3_2329,addr_selector3_2330,addr_selector3_2331,addr_selector3_2332,addr_selector3_2333,addr_selector3_2334,addr_selector3_2335,addr_selector3_2336,addr_selector3_2337,addr_selector3_2338,addr_selector3_2339,addr_selector3_2340,addr_selector3_2341,addr_selector3_2342,addr_selector3_2343,addr_selector3_2344,addr_selector3_2345,addr_selector3_2346,addr_selector3_2347,addr_selector3_2348,addr_selector3_2349,addr_selector3_2350,addr_selector3_2351,addr_selector3_2352,addr_selector3_2353,addr_selector3_2354,addr_selector3_2355,addr_selector3_2356,addr_selector3_2357,addr_selector3_2358,addr_selector3_2359,addr_selector3_2360,addr_selector3_2361,addr_selector3_2362,addr_selector3_2363,addr_selector3_2364,addr_selector3_2365,addr_selector3_2366,addr_selector3_2367,addr_selector3_2368,addr_selector3_2369,addr_selector3_2370,addr_selector3_2371,addr_selector3_2372,addr_selector3_2373,addr_selector3_2374,addr_selector3_2375,addr_selector3_2376,addr_selector3_2377,addr_selector3_2378,addr_selector3_2379,addr_selector3_2380,addr_selector3_2381,addr_selector3_2382,addr_selector3_2383,addr_selector3_2384,addr_selector3_2385,addr_selector3_2386,addr_selector3_2387,addr_selector3_2388,addr_selector3_2389,addr_selector3_2390,addr_selector3_2391,addr_selector3_2392,addr_selector3_2393,addr_selector3_2394,addr_selector3_2395,addr_selector3_2396,addr_selector3_2397,addr_selector3_2398,addr_selector3_2399,addr_selector3_2400,addr_selector3_2401,addr_selector3_2402,addr_selector3_2403,addr_selector3_2404,addr_selector3_2405,addr_selector3_2406,addr_selector3_2407,addr_selector3_2408,addr_selector3_2409,addr_selector3_2410,addr_selector3_2411,addr_selector3_2412,addr_selector3_2413,addr_selector3_2414,addr_selector3_2415,addr_selector3_2416,addr_selector3_2417,addr_selector3_2418,addr_selector3_2419,addr_selector3_2420,addr_selector3_2421,addr_selector3_2422,addr_selector3_2423,addr_selector3_2424,addr_selector3_2425,addr_selector3_2426,addr_selector3_2427,addr_selector3_2428,addr_selector3_2429,addr_selector3_2430,addr_selector3_2431,addr_selector3_2432,addr_selector3_2433,addr_selector3_2434,addr_selector3_2435,addr_selector3_2436,addr_selector3_2437,addr_selector3_2438,addr_selector3_2439,addr_selector3_2440,addr_selector3_2441,addr_selector3_2442,addr_selector3_2443,addr_selector3_2444,addr_selector3_2445,addr_selector3_2446,addr_selector3_2447,addr_selector3_2448,addr_selector3_2449,addr_selector3_2450,addr_selector3_2451,addr_selector3_2452,addr_selector3_2453,addr_selector3_2454,addr_selector3_2455,addr_selector3_2456,addr_selector3_2457,addr_selector3_2458,addr_selector3_2459,addr_selector3_2460,addr_selector3_2461,addr_selector3_2462,addr_selector3_2463,addr_selector3_2464,addr_selector3_2465,addr_selector3_2466,addr_selector3_2467,addr_selector3_2468,addr_selector3_2469,addr_selector3_2470,addr_selector3_2471,addr_selector3_2472,addr_selector3_2473,addr_selector3_2474,addr_selector3_2475,addr_selector3_2476,addr_selector3_2477,addr_selector3_2478,addr_selector3_2479,addr_selector3_2480,addr_selector3_2481,addr_selector3_2482,addr_selector3_2483,addr_selector3_2484,addr_selector3_2485,addr_selector3_2486,addr_selector3_2487,addr_selector3_2488,addr_selector3_2489,addr_selector3_2490,addr_selector3_2491,addr_selector3_2492,addr_selector3_2493,addr_selector3_2494,addr_selector3_2495,addr_selector3_2496,addr_selector3_2497,addr_selector3_2498,addr_selector3_2499,addr_selector3_2500,addr_selector3_2501,addr_selector3_2502,addr_selector3_2503,addr_selector3_2504,addr_selector3_2505,addr_selector3_2506,addr_selector3_2507,addr_selector3_2508,addr_selector3_2509,addr_selector3_2510,addr_selector3_2511,addr_selector3_2512,addr_selector3_2513,addr_selector3_2514,addr_selector3_2515,addr_selector3_2516,addr_selector3_2517,addr_selector3_2518,addr_selector3_2519,addr_selector3_2520,addr_selector3_2521,addr_selector3_2522,addr_selector3_2523,addr_selector3_2524,addr_selector3_2525,addr_selector3_2526,addr_selector3_2527,addr_selector3_2528,addr_selector3_2529,addr_selector3_2530,addr_selector3_2531,addr_selector3_2532,addr_selector3_2533,addr_selector3_2534,addr_selector3_2535,addr_selector3_2536,addr_selector3_2537,addr_selector3_2538,addr_selector3_2539,addr_selector3_2540,addr_selector3_2541,addr_selector3_2542,addr_selector3_2543,addr_selector3_2544,addr_selector3_2545,addr_selector3_2546,addr_selector3_2547,addr_selector3_2548,addr_selector3_2549,addr_selector3_2550,addr_selector3_2551,addr_selector3_2552,addr_selector3_2553,addr_selector3_2554,addr_selector3_2555,addr_selector3_2556,addr_selector3_2557,addr_selector3_2558,addr_selector3_2559,addr_selector3_2560,addr_selector3_2561,addr_selector3_2562,addr_selector3_2563,addr_selector3_2564,addr_selector3_2565,addr_selector3_2566,addr_selector3_2567,addr_selector3_2568,addr_selector3_2569,addr_selector3_2570,addr_selector3_2571,addr_selector3_2572,addr_selector3_2573,addr_selector3_2574,addr_selector3_2575,addr_selector3_2576,addr_selector3_2577,addr_selector3_2578,addr_selector3_2579,addr_selector3_2580,addr_selector3_2581,addr_selector3_2582,addr_selector3_2583,addr_selector3_2584,addr_selector3_2585,addr_selector3_2586,addr_selector3_2587,addr_selector3_2588,addr_selector3_2589,addr_selector3_2590,addr_selector3_2591,addr_selector3_2592,addr_selector3_2593,addr_selector3_2594,addr_selector3_2595,addr_selector3_2596,addr_selector3_2597,addr_selector3_2598,addr_selector3_2599,addr_selector3_2600,addr_selector3_2601,addr_selector3_2602,addr_selector3_2603,addr_selector3_2604,addr_selector3_2605,addr_selector3_2606,addr_selector3_2607,addr_selector3_2608,addr_selector3_2609,addr_selector3_2610,addr_selector3_2611,addr_selector3_2612,addr_selector3_2613,addr_selector3_2614,addr_selector3_2615,addr_selector3_2616,addr_selector3_2617,addr_selector3_2618,addr_selector3_2619,addr_selector3_2620,addr_selector3_2621,addr_selector3_2622,addr_selector3_2623,addr_selector3_2624,addr_selector3_2625,addr_selector3_2626,addr_selector3_2627,addr_selector3_2628,addr_selector3_2629,addr_selector3_2630,addr_selector3_2631,addr_selector3_2632,addr_selector3_2633,addr_selector3_2634,addr_selector3_2635,addr_selector3_2636,addr_selector3_2637,addr_selector3_2638,addr_selector3_2639,addr_selector3_2640,addr_selector3_2641,addr_selector3_2642,addr_selector3_2643,addr_selector3_2644,addr_selector3_2645,addr_selector3_2646,addr_selector3_2647,addr_selector3_2648,addr_selector3_2649,addr_selector3_2650,addr_selector3_2651,addr_selector3_2652,addr_selector3_2653,addr_selector3_2654,addr_selector3_2655,addr_selector3_2656,addr_selector3_2657,addr_selector3_2658,addr_selector3_2659,addr_selector3_2660,addr_selector3_2661,addr_selector3_2662,addr_selector3_2663,addr_selector3_2664,addr_selector3_2665,addr_selector3_2666,addr_selector3_2667,addr_selector3_2668,addr_selector3_2669,addr_selector3_2670,addr_selector3_2671,addr_selector3_2672,addr_selector3_2673,addr_selector3_2674,addr_selector3_2675,addr_selector3_2676,addr_selector3_2677,addr_selector3_2678,addr_selector3_2679,addr_selector3_2680,addr_selector3_2681,addr_selector3_2682,addr_selector3_2683,addr_selector3_2684,addr_selector3_2685,addr_selector3_2686,addr_selector3_2687,addr_selector3_2688,addr_selector3_2689,addr_selector3_2690,addr_selector3_2691,addr_selector3_2692,addr_selector3_2693,addr_selector3_2694,addr_selector3_2695,addr_selector3_2696,addr_selector3_2697,addr_selector3_2698,addr_selector3_2699,addr_selector3_2700,addr_selector3_2701,addr_selector3_2702,addr_selector3_2703,addr_selector3_2704,addr_selector3_2705,addr_selector3_2706,addr_selector3_2707,addr_selector3_2708,addr_selector3_2709,addr_selector3_2710,addr_selector3_2711,addr_selector3_2712,addr_selector3_2713,addr_selector3_2714,addr_selector3_2715,addr_selector3_2716,addr_selector3_2717,addr_selector3_2718,addr_selector3_2719,addr_selector3_2720,addr_selector3_2721,addr_selector3_2722,addr_selector3_2723,addr_selector3_2724,addr_selector3_2725,addr_selector3_2726,addr_selector3_2727,addr_selector3_2728,addr_selector3_2729,addr_selector3_2730,addr_selector3_2731,addr_selector3_2732,addr_selector3_2733,addr_selector3_2734,addr_selector3_2735,addr_selector3_2736,addr_selector3_2737,addr_selector3_2738,addr_selector3_2739,addr_selector3_2740,addr_selector3_2741,addr_selector3_2742,addr_selector3_2743,addr_selector3_2744,addr_selector3_2745,addr_selector3_2746,addr_selector3_2747,addr_selector3_2748,addr_selector3_2749,addr_selector3_2750,addr_selector3_2751,addr_selector3_2752,addr_selector3_2753,addr_selector3_2754,addr_selector3_2755,addr_selector3_2756,addr_selector3_2757,addr_selector3_2758,addr_selector3_2759,addr_selector3_2760,addr_selector3_2761,addr_selector3_2762,addr_selector3_2763,addr_selector3_2764,addr_selector3_2765,addr_selector3_2766,addr_selector3_2767,addr_selector3_2768,addr_selector3_2769,addr_selector3_2770,addr_selector3_2771,addr_selector3_2772,addr_selector3_2773,addr_selector3_2774,addr_selector3_2775,addr_selector3_2776,addr_selector3_2777,addr_selector3_2778,addr_selector3_2779,addr_selector3_2780,addr_selector3_2781,addr_selector3_2782,addr_selector3_2783,addr_selector3_2784,addr_selector3_2785,addr_selector3_2786,addr_selector3_2787,addr_selector3_2788,addr_selector3_2789,addr_selector3_2790,addr_selector3_2791,addr_selector3_2792,addr_selector3_2793,addr_selector3_2794,addr_selector3_2795,addr_selector3_2796,addr_selector3_2797,addr_selector3_2798,addr_selector3_2799,addr_selector3_2800,addr_selector3_2801,addr_selector3_2802,addr_selector3_2803,addr_selector3_2804,addr_selector3_2805,addr_selector3_2806,addr_selector3_2807,addr_selector3_2808,addr_selector3_2809,addr_selector3_2810,addr_selector3_2811,addr_selector3_2812,addr_selector3_2813,addr_selector3_2814,addr_selector3_2815,addr_selector3_2816,addr_selector3_2817,addr_selector3_2818,addr_selector3_2819,addr_selector3_2820,addr_selector3_2821,addr_selector3_2822,addr_selector3_2823,addr_selector3_2824,addr_selector3_2825,addr_selector3_2826,addr_selector3_2827,addr_selector3_2828,addr_selector3_2829,addr_selector3_2830,addr_selector3_2831,addr_selector3_2832,addr_selector3_2833,addr_selector3_2834,addr_selector3_2835,addr_selector3_2836,addr_selector3_2837,addr_selector3_2838,addr_selector3_2839,addr_selector3_2840,addr_selector3_2841,addr_selector3_2842,addr_selector3_2843,addr_selector3_2844,addr_selector3_2845,addr_selector3_2846,addr_selector3_2847,addr_selector3_2848,addr_selector3_2849,addr_selector3_2850,addr_selector3_2851,addr_selector3_2852,addr_selector3_2853,addr_selector3_2854,addr_selector3_2855,addr_selector3_2856,addr_selector3_2857,addr_selector3_2858,addr_selector3_2859,addr_selector3_2860,addr_selector3_2861,addr_selector3_2862,addr_selector3_2863,addr_selector3_2864,addr_selector3_2865,addr_selector3_2866,addr_selector3_2867,addr_selector3_2868,addr_selector3_2869,addr_selector3_2870,addr_selector3_2871,addr_selector3_2872,addr_selector3_2873,addr_selector3_2874,addr_selector3_2875,addr_selector3_2876,addr_selector3_2877,addr_selector3_2878,addr_selector3_2879,addr_selector3_2880,addr_selector3_2881,addr_selector3_2882,addr_selector3_2883,addr_selector3_2884,addr_selector3_2885,addr_selector3_2886,addr_selector3_2887,addr_selector3_2888,addr_selector3_2889,addr_selector3_2890,addr_selector3_2891,addr_selector3_2892,addr_selector3_2893,addr_selector3_2894,addr_selector3_2895,addr_selector3_2896,addr_selector3_2897,addr_selector3_2898,addr_selector3_2899,addr_selector3_2900,addr_selector3_2901,addr_selector3_2902,addr_selector3_2903,addr_selector3_2904,addr_selector3_2905,addr_selector3_2906,addr_selector3_2907,addr_selector3_2908,addr_selector3_2909,addr_selector3_2910,addr_selector3_2911,addr_selector3_2912,addr_selector3_2913,addr_selector3_2914,addr_selector3_2915,addr_selector3_2916,addr_selector3_2917,addr_selector3_2918,addr_selector3_2919,addr_selector3_2920,addr_selector3_2921,addr_selector3_2922,addr_selector3_2923,addr_selector3_2924,addr_selector3_2925,addr_selector3_2926,addr_selector3_2927,addr_selector3_2928,addr_selector3_2929,addr_selector3_2930,addr_selector3_2931,addr_selector3_2932,addr_selector3_2933,addr_selector3_2934,addr_selector3_2935,addr_selector3_2936,addr_selector3_2937,addr_selector3_2938,addr_selector3_2939,addr_selector3_2940,addr_selector3_2941,addr_selector3_2942,addr_selector3_2943,addr_selector3_2944,addr_selector3_2945,addr_selector3_2946,addr_selector3_2947,addr_selector3_2948,addr_selector3_2949,addr_selector3_2950,addr_selector3_2951,addr_selector3_2952,addr_selector3_2953,addr_selector3_2954,addr_selector3_2955,addr_selector3_2956,addr_selector3_2957,addr_selector3_2958,addr_selector3_2959,addr_selector3_2960,addr_selector3_2961,addr_selector3_2962,addr_selector3_2963,addr_selector3_2964,addr_selector3_2965,addr_selector3_2966,addr_selector3_2967,addr_selector3_2968,addr_selector3_2969,addr_selector3_2970,addr_selector3_2971,addr_selector3_2972,addr_selector3_2973,addr_selector3_2974,addr_selector3_2975,addr_selector3_2976,addr_selector3_2977,addr_selector3_2978,addr_selector3_2979,addr_selector3_2980,addr_selector3_2981,addr_selector3_2982,addr_selector3_2983,addr_selector3_2984,addr_selector3_2985,addr_selector3_2986,addr_selector3_2987,addr_selector3_2988,addr_selector3_2989,addr_selector3_2990,addr_selector3_2991,addr_selector3_2992,addr_selector3_2993,addr_selector3_2994,addr_selector3_2995,addr_selector3_2996,addr_selector3_2997,addr_selector3_2998,addr_selector3_2999,addr_selector3_3000,addr_selector3_3001,addr_selector3_3002,addr_selector3_3003,addr_selector3_3004,addr_selector3_3005,addr_selector3_3006,addr_selector3_3007,addr_selector3_3008,addr_selector3_3009,addr_selector3_3010,addr_selector3_3011,addr_selector3_3012,addr_selector3_3013,addr_selector3_3014,addr_selector3_3015,addr_selector3_3016,addr_selector3_3017,addr_selector3_3018,addr_selector3_3019,addr_selector3_3020,addr_selector3_3021,addr_selector3_3022,addr_selector3_3023,addr_selector3_3024,addr_selector3_3025,addr_selector3_3026,addr_selector3_3027,addr_selector3_3028,addr_selector3_3029,addr_selector3_3030,addr_selector3_3031,addr_selector3_3032,addr_selector3_3033,addr_selector3_3034,addr_selector3_3035,addr_selector3_3036,addr_selector3_3037,addr_selector3_3038,addr_selector3_3039,addr_selector3_3040,addr_selector3_3041,addr_selector3_3042,addr_selector3_3043,addr_selector3_3044,addr_selector3_3045,addr_selector3_3046,addr_selector3_3047,addr_selector3_3048,addr_selector3_3049,addr_selector3_3050,addr_selector3_3051,addr_selector3_3052,addr_selector3_3053,addr_selector3_3054,addr_selector3_3055,addr_selector3_3056,addr_selector3_3057,addr_selector3_3058,addr_selector3_3059,addr_selector3_3060,addr_selector3_3061,addr_selector3_3062,addr_selector3_3063,addr_selector3_3064,addr_selector3_3065,addr_selector3_3066,addr_selector3_3067,addr_selector3_3068,addr_selector3_3069,addr_selector3_3070,addr_selector3_3071,addr_selector3_3072,addr_selector3_3073,addr_selector3_3074,addr_selector3_3075,addr_selector3_3076,addr_selector3_3077,addr_selector3_3078,addr_selector3_3079,addr_selector3_3080,addr_selector3_3081,addr_selector3_3082,addr_selector3_3083,addr_selector3_3084,addr_selector3_3085,addr_selector3_3086,addr_selector3_3087,addr_selector3_3088,addr_selector3_3089,addr_selector3_3090,addr_selector3_3091,addr_selector3_3092,addr_selector3_3093,addr_selector3_3094,addr_selector3_3095,addr_selector3_3096,addr_selector3_3097,addr_selector3_3098,addr_selector3_3099,addr_selector3_3100,addr_selector3_3101,addr_selector3_3102,addr_selector3_3103,addr_selector3_3104,addr_selector3_3105,addr_selector3_3106,addr_selector3_3107,addr_selector3_3108,addr_selector3_3109,addr_selector3_3110,addr_selector3_3111,addr_selector3_3112,addr_selector3_3113,addr_selector3_3114,addr_selector3_3115,addr_selector3_3116,addr_selector3_3117,addr_selector3_3118,addr_selector3_3119,addr_selector3_3120,addr_selector3_3121,addr_selector3_3122,addr_selector3_3123,addr_selector3_3124,addr_selector3_3125,addr_selector3_3126,addr_selector3_3127,addr_selector3_3128,addr_selector3_3129,addr_selector3_3130,addr_selector3_3131,addr_selector3_3132,addr_selector3_3133,addr_selector3_3134,addr_selector3_3135,addr_selector3_3136,addr_selector3_3137,addr_selector3_3138,addr_selector3_3139,addr_selector3_3140,addr_selector3_3141,addr_selector3_3142,addr_selector3_3143,addr_selector3_3144,addr_selector3_3145,addr_selector3_3146,addr_selector3_3147,addr_selector3_3148,addr_selector3_3149,addr_selector3_3150,addr_selector3_3151,addr_selector3_3152,addr_selector3_3153,addr_selector3_3154,addr_selector3_3155,addr_selector3_3156,addr_selector3_3157,addr_selector3_3158,addr_selector3_3159,addr_selector3_3160,addr_selector3_3161,addr_selector3_3162,addr_selector3_3163,addr_selector3_3164,addr_selector3_3165,addr_selector3_3166,addr_selector3_3167,addr_selector3_3168,addr_selector3_3169,addr_selector3_3170,addr_selector3_3171,addr_selector3_3172,addr_selector3_3173,addr_selector3_3174,addr_selector3_3175,addr_selector3_3176,addr_selector3_3177,addr_selector3_3178,addr_selector3_3179,addr_selector3_3180,addr_selector3_3181,addr_selector3_3182,addr_selector3_3183,addr_selector3_3184,addr_selector3_3185,addr_selector3_3186,addr_selector3_3187,addr_selector3_3188,addr_selector3_3189,addr_selector3_3190,addr_selector3_3191,addr_selector3_3192,addr_selector3_3193,addr_selector3_3194,addr_selector3_3195,addr_selector3_3196,addr_selector3_3197,addr_selector3_3198,addr_selector3_3199,addr_selector3_3200,addr_selector3_3201,addr_selector3_3202,addr_selector3_3203,addr_selector3_3204,addr_selector3_3205,addr_selector3_3206,addr_selector3_3207,addr_selector3_3208,addr_selector3_3209,addr_selector3_3210,addr_selector3_3211,addr_selector3_3212,addr_selector3_3213,addr_selector3_3214,addr_selector3_3215,addr_selector3_3216,addr_selector3_3217,addr_selector3_3218,addr_selector3_3219,addr_selector3_3220,addr_selector3_3221,addr_selector3_3222,addr_selector3_3223,addr_selector3_3224,addr_selector3_3225,addr_selector3_3226,addr_selector3_3227,addr_selector3_3228,addr_selector3_3229,addr_selector3_3230,addr_selector3_3231,addr_selector3_3232,addr_selector3_3233,addr_selector3_3234,addr_selector3_3235,addr_selector3_3236,addr_selector3_3237,addr_selector3_3238,addr_selector3_3239,addr_selector3_3240,addr_selector3_3241,addr_selector3_3242,addr_selector3_3243,addr_selector3_3244,addr_selector3_3245,addr_selector3_3246,addr_selector3_3247,addr_selector3_3248,addr_selector3_3249,addr_selector3_3250,addr_selector3_3251,addr_selector3_3252,addr_selector3_3253,addr_selector3_3254,addr_selector3_3255,addr_selector3_3256,addr_selector3_3257,addr_selector3_3258,addr_selector3_3259,addr_selector3_3260,addr_selector3_3261,addr_selector3_3262,addr_selector3_3263,addr_selector3_3264,addr_selector3_3265,addr_selector3_3266,addr_selector3_3267,addr_selector3_3268,addr_selector3_3269,addr_selector3_3270,addr_selector3_3271,addr_selector3_3272,addr_selector3_3273,addr_selector3_3274,addr_selector3_3275,addr_selector3_3276,addr_selector3_3277,addr_selector3_3278,addr_selector3_3279,addr_selector3_3280,addr_selector3_3281,addr_selector3_3282,addr_selector3_3283,addr_selector3_3284,addr_selector3_3285,addr_selector3_3286,addr_selector3_3287,addr_selector3_3288,addr_selector3_3289,addr_selector3_3290,addr_selector3_3291,addr_selector3_3292,addr_selector3_3293,addr_selector3_3294,addr_selector3_3295,addr_selector3_3296,addr_selector3_3297,addr_selector3_3298,addr_selector3_3299,addr_selector3_3300,addr_selector3_3301,addr_selector3_3302,addr_selector3_3303,addr_selector3_3304,addr_selector3_3305,addr_selector3_3306,addr_selector3_3307,addr_selector3_3308,addr_selector3_3309,addr_selector3_3310,addr_selector3_3311,addr_selector3_3312,addr_selector3_3313,addr_selector3_3314,addr_selector3_3315,addr_selector3_3316,addr_selector3_3317,addr_selector3_3318,addr_selector3_3319,addr_selector3_3320,addr_selector3_3321,addr_selector3_3322,addr_selector3_3323,addr_selector3_3324,addr_selector3_3325,addr_selector3_3326,addr_selector3_3327,addr_selector3_3328,addr_selector3_3329,addr_selector3_3330,addr_selector3_3331,addr_selector3_3332,addr_selector3_3333,addr_selector3_3334,addr_selector3_3335,addr_selector3_3336,addr_selector3_3337,addr_selector3_3338,addr_selector3_3339,addr_selector3_3340,addr_selector3_3341,addr_selector3_3342,addr_selector3_3343,addr_selector3_3344,addr_selector3_3345,addr_selector3_3346,addr_selector3_3347,addr_selector3_3348,addr_selector3_3349,addr_selector3_3350,addr_selector3_3351,addr_selector3_3352,addr_selector3_3353,addr_selector3_3354,addr_selector3_3355,addr_selector3_3356,addr_selector3_3357,addr_selector3_3358,addr_selector3_3359,addr_selector3_3360,addr_selector3_3361,addr_selector3_3362,addr_selector3_3363,addr_selector3_3364,addr_selector3_3365,addr_selector3_3366,addr_selector3_3367,addr_selector3_3368,addr_selector3_3369,addr_selector3_3370,addr_selector3_3371,addr_selector3_3372,addr_selector3_3373,addr_selector3_3374,addr_selector3_3375,addr_selector3_3376,addr_selector3_3377,addr_selector3_3378,addr_selector3_3379,addr_selector3_3380,addr_selector3_3381,addr_selector3_3382,addr_selector3_3383,addr_selector3_3384,addr_selector3_3385,addr_selector3_3386,addr_selector3_3387,addr_selector3_3388,addr_selector3_3389,addr_selector3_3390,addr_selector3_3391,addr_selector3_3392,addr_selector3_3393,addr_selector3_3394,addr_selector3_3395,addr_selector3_3396,addr_selector3_3397,addr_selector3_3398,addr_selector3_3399,addr_selector3_3400,addr_selector3_3401,addr_selector3_3402,addr_selector3_3403,addr_selector3_3404,addr_selector3_3405,addr_selector3_3406,addr_selector3_3407,addr_selector3_3408,addr_selector3_3409,addr_selector3_3410,addr_selector3_3411,addr_selector3_3412,addr_selector3_3413,addr_selector3_3414,addr_selector3_3415,addr_selector3_3416,addr_selector3_3417,addr_selector3_3418,addr_selector3_3419,addr_selector3_3420,addr_selector3_3421,addr_selector3_3422,addr_selector3_3423,addr_selector3_3424,addr_selector3_3425,addr_selector3_3426,addr_selector3_3427,addr_selector3_3428,addr_selector3_3429,addr_selector3_3430,addr_selector3_3431,addr_selector3_3432,addr_selector3_3433,addr_selector3_3434,addr_selector3_3435,addr_selector3_3436,addr_selector3_3437,addr_selector3_3438,addr_selector3_3439,addr_selector3_3440,addr_selector3_3441,addr_selector3_3442,addr_selector3_3443,addr_selector3_3444,addr_selector3_3445,addr_selector3_3446,addr_selector3_3447,addr_selector3_3448,addr_selector3_3449,addr_selector3_3450,addr_selector3_3451,addr_selector3_3452,addr_selector3_3453,addr_selector3_3454,addr_selector3_3455,addr_selector3_3456,addr_selector3_3457,addr_selector3_3458,addr_selector3_3459,addr_selector3_3460,addr_selector3_3461,addr_selector3_3462,addr_selector3_3463,addr_selector3_3464,addr_selector3_3465,addr_selector3_3466,addr_selector3_3467,addr_selector3_3468,addr_selector3_3469,addr_selector3_3470,addr_selector3_3471,addr_selector3_3472,addr_selector3_3473,addr_selector3_3474,addr_selector3_3475,addr_selector3_3476,addr_selector3_3477,addr_selector3_3478,addr_selector3_3479,addr_selector3_3480,addr_selector3_3481,addr_selector3_3482,addr_selector3_3483,addr_selector3_3484,addr_selector3_3485,addr_selector3_3486,addr_selector3_3487,addr_selector3_3488,addr_selector3_3489,addr_selector3_3490,addr_selector3_3491,addr_selector3_3492,addr_selector3_3493,addr_selector3_3494,addr_selector3_3495,addr_selector3_3496,addr_selector3_3497,addr_selector3_3498,addr_selector3_3499,addr_selector3_3500,addr_selector3_3501,addr_selector3_3502,addr_selector3_3503,addr_selector3_3504,addr_selector3_3505,addr_selector3_3506,addr_selector3_3507,addr_selector3_3508,addr_selector3_3509,addr_selector3_3510,addr_selector3_3511,addr_selector3_3512,addr_selector3_3513,addr_selector3_3514,addr_selector3_3515,addr_selector3_3516,addr_selector3_3517,addr_selector3_3518,addr_selector3_3519,addr_selector3_3520,addr_selector3_3521,addr_selector3_3522,addr_selector3_3523,addr_selector3_3524,addr_selector3_3525,addr_selector3_3526,addr_selector3_3527,addr_selector3_3528,addr_selector3_3529,addr_selector3_3530,addr_selector3_3531,addr_selector3_3532,addr_selector3_3533,addr_selector3_3534,addr_selector3_3535,addr_selector3_3536,addr_selector3_3537,addr_selector3_3538,addr_selector3_3539,addr_selector3_3540,addr_selector3_3541,addr_selector3_3542,addr_selector3_3543,addr_selector3_3544,addr_selector3_3545,addr_selector3_3546,addr_selector3_3547,addr_selector3_3548,addr_selector3_3549,addr_selector3_3550,addr_selector3_3551,addr_selector3_3552,addr_selector3_3553,addr_selector3_3554,addr_selector3_3555,addr_selector3_3556,addr_selector3_3557,addr_selector3_3558,addr_selector3_3559,addr_selector3_3560,addr_selector3_3561,addr_selector3_3562,addr_selector3_3563,addr_selector3_3564,addr_selector3_3565,addr_selector3_3566,addr_selector3_3567,addr_selector3_3568,addr_selector3_3569,addr_selector3_3570,addr_selector3_3571,addr_selector3_3572,addr_selector3_3573,addr_selector3_3574,addr_selector3_3575,addr_selector3_3576,addr_selector3_3577,addr_selector3_3578,addr_selector3_3579,addr_selector3_3580,addr_selector3_3581,addr_selector3_3582,addr_selector3_3583,addr_selector3_3584,addr_selector3_3585,addr_selector3_3586,addr_selector3_3587,addr_selector3_3588,addr_selector3_3589,addr_selector3_3590,addr_selector3_3591,addr_selector3_3592,addr_selector3_3593,addr_selector3_3594,addr_selector3_3595,addr_selector3_3596,addr_selector3_3597,addr_selector3_3598,addr_selector3_3599,addr_selector3_3600,addr_selector3_3601,addr_selector3_3602,addr_selector3_3603,addr_selector3_3604,addr_selector3_3605,addr_selector3_3606,addr_selector3_3607,addr_selector3_3608,addr_selector3_3609,addr_selector3_3610,addr_selector3_3611,addr_selector3_3612,addr_selector3_3613,addr_selector3_3614,addr_selector3_3615,addr_selector3_3616,addr_selector3_3617,addr_selector3_3618,addr_selector3_3619,addr_selector3_3620,addr_selector3_3621,addr_selector3_3622,addr_selector3_3623,addr_selector3_3624,addr_selector3_3625,addr_selector3_3626,addr_selector3_3627,addr_selector3_3628,addr_selector3_3629,addr_selector3_3630,addr_selector3_3631,addr_selector3_3632,addr_selector3_3633,addr_selector3_3634,addr_selector3_3635,addr_selector3_3636,addr_selector3_3637,addr_selector3_3638,addr_selector3_3639,addr_selector3_3640,addr_selector3_3641,addr_selector3_3642,addr_selector3_3643,addr_selector3_3644,addr_selector3_3645,addr_selector3_3646,addr_selector3_3647,addr_selector3_3648,addr_selector3_3649,addr_selector3_3650,addr_selector3_3651,addr_selector3_3652,addr_selector3_3653,addr_selector3_3654,addr_selector3_3655,addr_selector3_3656,addr_selector3_3657,addr_selector3_3658,addr_selector3_3659,addr_selector3_3660,addr_selector3_3661,addr_selector3_3662,addr_selector3_3663,addr_selector3_3664,addr_selector3_3665,addr_selector3_3666,addr_selector3_3667,addr_selector3_3668,addr_selector3_3669,addr_selector3_3670,addr_selector3_3671,addr_selector3_3672,addr_selector3_3673,addr_selector3_3674,addr_selector3_3675,addr_selector3_3676,addr_selector3_3677,addr_selector3_3678,addr_selector3_3679,addr_selector3_3680,addr_selector3_3681,addr_selector3_3682,addr_selector3_3683,addr_selector3_3684,addr_selector3_3685,addr_selector3_3686,addr_selector3_3687,addr_selector3_3688,addr_selector3_3689,addr_selector3_3690,addr_selector3_3691,addr_selector3_3692,addr_selector3_3693,addr_selector3_3694,addr_selector3_3695,addr_selector3_3696,addr_selector3_3697,addr_selector3_3698,addr_selector3_3699,addr_selector3_3700,addr_selector3_3701,addr_selector3_3702,addr_selector3_3703,addr_selector3_3704,addr_selector3_3705,addr_selector3_3706,addr_selector3_3707,addr_selector3_3708,addr_selector3_3709,addr_selector3_3710,addr_selector3_3711,addr_selector3_3712,addr_selector3_3713,addr_selector3_3714,addr_selector3_3715,addr_selector3_3716,addr_selector3_3717,addr_selector3_3718,addr_selector3_3719,addr_selector3_3720,addr_selector3_3721,addr_selector3_3722,addr_selector3_3723,addr_selector3_3724,addr_selector3_3725,addr_selector3_3726,addr_selector3_3727,addr_selector3_3728,addr_selector3_3729,addr_selector3_3730,addr_selector3_3731,addr_selector3_3732,addr_selector3_3733,addr_selector3_3734,addr_selector3_3735,addr_selector3_3736,addr_selector3_3737,addr_selector3_3738,addr_selector3_3739,addr_selector3_3740,addr_selector3_3741,addr_selector3_3742,addr_selector3_3743,addr_selector3_3744,addr_selector3_3745,addr_selector3_3746,addr_selector3_3747,addr_selector3_3748,addr_selector3_3749,addr_selector3_3750,addr_selector3_3751,addr_selector3_3752,addr_selector3_3753,addr_selector3_3754,addr_selector3_3755,addr_selector3_3756,addr_selector3_3757,addr_selector3_3758,addr_selector3_3759,addr_selector3_3760,addr_selector3_3761,addr_selector3_3762,addr_selector3_3763,addr_selector3_3764,addr_selector3_3765,addr_selector3_3766,addr_selector3_3767,addr_selector3_3768,addr_selector3_3769,addr_selector3_3770,addr_selector3_3771,addr_selector3_3772,addr_selector3_3773,addr_selector3_3774,addr_selector3_3775,addr_selector3_3776,addr_selector3_3777,addr_selector3_3778,addr_selector3_3779,addr_selector3_3780,addr_selector3_3781,addr_selector3_3782,addr_selector3_3783,addr_selector3_3784,addr_selector3_3785,addr_selector3_3786,addr_selector3_3787,addr_selector3_3788,addr_selector3_3789,addr_selector3_3790,addr_selector3_3791,addr_selector3_3792,addr_selector3_3793,addr_selector3_3794,addr_selector3_3795,addr_selector3_3796,addr_selector3_3797,addr_selector3_3798,addr_selector3_3799,addr_selector3_3800,addr_selector3_3801,addr_selector3_3802,addr_selector3_3803,addr_selector3_3804,addr_selector3_3805,addr_selector3_3806,addr_selector3_3807,addr_selector3_3808,addr_selector3_3809,addr_selector3_3810,addr_selector3_3811,addr_selector3_3812,addr_selector3_3813,addr_selector3_3814,addr_selector3_3815,addr_selector3_3816,addr_selector3_3817,addr_selector3_3818,addr_selector3_3819,addr_selector3_3820,addr_selector3_3821,addr_selector3_3822,addr_selector3_3823,addr_selector3_3824,addr_selector3_3825,addr_selector3_3826,addr_selector3_3827,addr_selector3_3828,addr_selector3_3829,addr_selector3_3830,addr_selector3_3831,addr_selector3_3832,addr_selector3_3833,addr_selector3_3834,addr_selector3_3835,addr_selector3_3836,addr_selector3_3837,addr_selector3_3838,addr_selector3_3839,addr_selector3_3840,addr_selector3_3841,addr_selector3_3842,addr_selector3_3843,addr_selector3_3844,addr_selector3_3845,addr_selector3_3846,addr_selector3_3847,addr_selector3_3848,addr_selector3_3849,addr_selector3_3850,addr_selector3_3851,addr_selector3_3852,addr_selector3_3853,addr_selector3_3854,addr_selector3_3855,addr_selector3_3856,addr_selector3_3857,addr_selector3_3858,addr_selector3_3859,addr_selector3_3860,addr_selector3_3861,addr_selector3_3862,addr_selector3_3863,addr_selector3_3864,addr_selector3_3865,addr_selector3_3866,addr_selector3_3867,addr_selector3_3868,addr_selector3_3869,addr_selector3_3870,addr_selector3_3871,addr_selector3_3872,addr_selector3_3873,addr_selector3_3874,addr_selector3_3875,addr_selector3_3876,addr_selector3_3877,addr_selector3_3878,addr_selector3_3879,addr_selector3_3880,addr_selector3_3881,addr_selector3_3882,addr_selector3_3883,addr_selector3_3884,addr_selector3_3885,addr_selector3_3886,addr_selector3_3887,addr_selector3_3888,addr_selector3_3889,addr_selector3_3890,addr_selector3_3891,addr_selector3_3892,addr_selector3_3893,addr_selector3_3894,addr_selector3_3895,addr_selector3_3896,addr_selector3_3897,addr_selector3_3898,addr_selector3_3899,addr_selector3_3900,addr_selector3_3901,addr_selector3_3902,addr_selector3_3903,addr_selector3_3904,addr_selector3_3905,addr_selector3_3906,addr_selector3_3907,addr_selector3_3908,addr_selector3_3909,addr_selector3_3910,addr_selector3_3911,addr_selector3_3912,addr_selector3_3913,addr_selector3_3914,addr_selector3_3915,addr_selector3_3916,addr_selector3_3917,addr_selector3_3918,addr_selector3_3919,addr_selector3_3920,addr_selector3_3921,addr_selector3_3922,addr_selector3_3923,addr_selector3_3924,addr_selector3_3925,addr_selector3_3926,addr_selector3_3927,addr_selector3_3928,addr_selector3_3929,addr_selector3_3930,addr_selector3_3931,addr_selector3_3932,addr_selector3_3933,addr_selector3_3934,addr_selector3_3935,addr_selector3_3936,addr_selector3_3937,addr_selector3_3938,addr_selector3_3939,addr_selector3_3940,addr_selector3_3941,addr_selector3_3942,addr_selector3_3943,addr_selector3_3944,addr_selector3_3945,addr_selector3_3946,addr_selector3_3947,addr_selector3_3948,addr_selector3_3949,addr_selector3_3950,addr_selector3_3951,addr_selector3_3952,addr_selector3_3953,addr_selector3_3954,addr_selector3_3955,addr_selector3_3956,addr_selector3_3957,addr_selector3_3958,addr_selector3_3959,addr_selector3_3960,addr_selector3_3961,addr_selector3_3962,addr_selector3_3963,addr_selector3_3964,addr_selector3_3965,addr_selector3_3966,addr_selector3_3967,addr_selector3_3968,addr_selector3_3969,addr_selector3_3970,addr_selector3_3971,addr_selector3_3972,addr_selector3_3973,addr_selector3_3974,addr_selector3_3975,addr_selector3_3976,addr_selector3_3977,addr_selector3_3978,addr_selector3_3979,addr_selector3_3980,addr_selector3_3981,addr_selector3_3982,addr_selector3_3983,addr_selector3_3984,addr_selector3_3985,addr_selector3_3986,addr_selector3_3987,addr_selector3_3988,addr_selector3_3989,addr_selector3_3990,addr_selector3_3991,addr_selector3_3992,addr_selector3_3993,addr_selector3_3994,addr_selector3_3995,addr_selector3_3996,addr_selector3_3997,addr_selector3_3998,addr_selector3_3999,addr_selector3_4000,addr_selector3_4001,addr_selector3_4002,addr_selector3_4003,addr_selector3_4004,addr_selector3_4005,addr_selector3_4006,addr_selector3_4007,addr_selector3_4008,addr_selector3_4009,addr_selector3_4010,addr_selector3_4011,addr_selector3_4012,addr_selector3_4013,addr_selector3_4014,addr_selector3_4015,addr_selector3_4016,addr_selector3_4017,addr_selector3_4018,addr_selector3_4019,addr_selector3_4020,addr_selector3_4021,addr_selector3_4022,addr_selector3_4023,addr_selector3_4024,addr_selector3_4025,addr_selector3_4026,addr_selector3_4027,addr_selector3_4028,addr_selector3_4029,addr_selector3_4030,addr_selector3_4031,addr_selector3_4032,addr_selector3_4033,addr_selector3_4034,addr_selector3_4035,addr_selector3_4036,addr_selector3_4037,addr_selector3_4038,addr_selector3_4039,addr_selector3_4040,addr_selector3_4041,addr_selector3_4042,addr_selector3_4043,addr_selector3_4044,addr_selector3_4045,addr_selector3_4046,addr_selector3_4047,addr_selector3_4048,addr_selector3_4049,addr_selector3_4050,addr_selector3_4051,addr_selector3_4052,addr_selector3_4053,addr_selector3_4054,addr_selector3_4055,addr_selector3_4056,addr_selector3_4057,addr_selector3_4058,addr_selector3_4059,addr_selector3_4060,addr_selector3_4061,addr_selector3_4062,addr_selector3_4063,addr_selector3_4064,addr_selector3_4065,addr_selector3_4066,addr_selector3_4067,addr_selector3_4068,addr_selector3_4069,addr_selector3_4070,addr_selector3_4071,addr_selector3_4072,addr_selector3_4073,addr_selector3_4074,addr_selector3_4075,addr_selector3_4076,addr_selector3_4077,addr_selector3_4078,addr_selector3_4079,addr_selector3_4080,addr_selector3_4081,addr_selector3_4082,addr_selector3_4083,addr_selector3_4084,addr_selector3_4085,addr_selector3_4086,addr_selector3_4087,addr_selector3_4088,addr_selector3_4089,addr_selector3_4090,addr_selector3_4091,addr_selector3_4092,addr_selector3_4093,addr_selector3_4094,addr_selector3_4095};


endmodule
